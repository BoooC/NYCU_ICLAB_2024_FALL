// ##############################################################
//   You can modify by your own
//   You can modify by your own
//   You can modify by your own
// ##############################################################

module CHIP(
    // input signals
    clk,
    rst_n,
    in_valid, 
    in_valid2,
    
    image,
    template,
    image_size,
	action,
	
    // output signals
    out_valid,
    out_value
);


input            clk, rst_n, in_valid, in_valid2;
input     [7:0]  image;
input     [7:0]  template;
input     [1:0]  image_size;
input     [2:0]  action;

output           out_valid;
output           out_value;

//==================================================================
// reg & wire
//==================================================================
wire             C_clk;
wire             C_rst_n;
wire             C_in_valid;
wire             C_in_valid2;

wire     [7:0]   C_image;
wire     [7:0]   C_template;
wire     [1:0]   C_image_size;
wire     [2:0]   C_action;

wire             C_out_valid;
wire             C_out_value;

//==================================================================
// CORE
//==================================================================
TMIP CORE(
	// input signals
    .clk(C_clk),
    .rst_n(C_rst_n),
    .in_valid(C_in_valid), 
    .in_valid2(C_in_valid2),
    
    .image(C_image),
    .template(C_template),
    .image_size(C_image_size),
	.action(C_action),
	
    // output signals
    .out_valid(C_out_valid),
    .out_value(C_out_value)
);

//==================================================================
// INPUT PAD
// Syntax: XMD PAD_NAME ( .O(CORE_PORT_NAME), .I(CHIP_PORT_NAME), .PU(1'b0), .PD(1'b0), .SMT(1'b0));
//     Ex: XMD    I_CLK ( .O(C_clk),          .I(clk),            .PU(1'b0), .PD(1'b0), .SMT(1'b0));
//==================================================================
// You need to finish this part
XMD    I_CLK        ( .O(C_clk),            .I(clk),            .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_RST        ( .O(C_rst_n),          .I(rst_n),          .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IN_VALID   ( .O(C_in_valid),       .I(in_valid),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IN_VALID2  ( .O(C_in_valid2),      .I(in_valid2),      .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE0     ( .O(C_image[0]),       .I(image[0]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE1     ( .O(C_image[1]),       .I(image[1]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE2     ( .O(C_image[2]),       .I(image[2]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE3     ( .O(C_image[3]),       .I(image[3]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE4     ( .O(C_image[4]),       .I(image[4]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE5     ( .O(C_image[5]),       .I(image[5]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE6     ( .O(C_image[6]),       .I(image[6]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE7     ( .O(C_image[7]),       .I(image[7]),       .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE0  ( .O(C_template[0]),    .I(template[0]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE1  ( .O(C_template[1]),    .I(template[1]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE2  ( .O(C_template[2]),    .I(template[2]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE3  ( .O(C_template[3]),    .I(template[3]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE4  ( .O(C_template[4]),    .I(template[4]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE5  ( .O(C_template[5]),    .I(template[5]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE6  ( .O(C_template[6]),    .I(template[6]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_TEMPLATE7  ( .O(C_template[7]),    .I(template[7]),    .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE_SIZE0( .O(C_image_size[0]),  .I(image_size[0]),  .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_IMAGE_SIZE1( .O(C_image_size[1]),  .I(image_size[1]),  .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_ACTION0    ( .O(C_action[0]),      .I(action[0]),      .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_ACTION1    ( .O(C_action[1]),      .I(action[1]),      .PU(1'b0), .PD(1'b0), .SMT(1'b0));
XMD    I_ACTION2    ( .O(C_action[2]),      .I(action[2]),      .PU(1'b0), .PD(1'b0), .SMT(1'b0));

//==================================================================
// OUTPUT PAD
// Syntax: YA2GSD PAD_NAME (.I(CORE_PIN_NAME), .O(PAD_PIN_NAME), .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
//     Ex: YA2GSD  O_VALID (.I(C_out_valid),   .O(out_valid),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
//==================================================================
// You need to finish this part
YA2GSD  O_VALID (.I(C_out_valid),   .O(out_valid),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));
YA2GSD  O_VALUE (.I(C_out_value),   .O(out_value),    .E(1'b1), .E2(1'b1), .E4(1'b1), .E8(1'b0), .SR(1'b0));

//==================================================================
// I/O power 3.3V pads x? (DVDD + DGND)
// Syntax: VCC3IOD/GNDIOD PAD_NAME ();
//    Ex1: VCC3IOD        VDDP0 ();
//    Ex2: GNDIOD         GNDP0 ();
//==================================================================
// You need to finish this part
VCC3IOD     VDDP0 ();
GNDIOD      GNDP0 ();
VCC3IOD     VDDP1 ();
GNDIOD      GNDP1 ();
VCC3IOD     VDDP2 ();
GNDIOD      GNDP2 ();
// VCC3IOD     VDDP3 ();
// GNDIOD      GNDP3 ();

//==================================================================
// Core power 1.8V pads x? (VDD + GND)
// Syntax: VCCKD/GNDKD PAD_NAME ();
//    Ex1: VCCKD       VDDC0 ();
//    Ex2: GNDKD       GNDC0 ();
//==================================================================
// You need to finish this part
VCCKD       VDDC0 ();
GNDKD       GNDC0 ();
VCCKD       VDDC1 ();
GNDKD       GNDC1 ();
// VCCKD       VDDC2 ();
// GNDKD       GNDC2 ();
// VCCKD       VDDC3 ();
// GNDKD       GNDC3 ();

endmodule

/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Ultra(TM) in wire load mode
// Version   : T-2022.03
// Date      : Mon Dec  2 02:57:51 2024
/////////////////////////////////////////////////////////////


module TMIP ( clk, rst_n, in_valid, in_valid2, image, template, image_size, 
        action, out_valid, out_value );
  input [7:0] image;
  input [7:0] template;
  input [1:0] image_size;
  input [2:0] action;
  input clk, rst_n, in_valid, in_valid2;
  output out_valid, out_value;
  wire   SRAM_192_32_read_done, flip_flag, neg_flag, window_0__3__7_,
         window_0__3__6_, window_0__3__5_, window_0__3__4_, window_0__3__3_,
         window_0__3__2_, window_0__3__1_, window_0__3__0_, window_0__4__7_,
         window_0__4__6_, window_0__4__5_, window_0__4__4_, window_0__4__3_,
         window_0__4__2_, window_0__4__1_, window_0__4__0_, window_1__3__7_,
         window_1__3__6_, window_1__3__5_, window_1__3__4_, window_1__3__3_,
         window_1__3__2_, window_1__3__1_, window_1__3__0_, window_1__4__7_,
         window_1__4__6_, window_1__4__5_, window_1__4__4_, window_1__4__3_,
         window_1__4__2_, window_1__4__1_, window_1__4__0_, window_2__3__7_,
         window_2__3__6_, window_2__3__5_, window_2__3__4_, window_2__3__3_,
         window_2__3__2_, window_2__3__1_, window_2__3__0_, window_2__4__7_,
         window_2__4__6_, window_2__4__5_, window_2__4__4_, window_2__4__3_,
         window_2__4__2_, window_2__4__1_, window_2__4__0_, action_reg_0__1_,
         action_reg_0__0_, action_reg_1__2_, action_reg_1__1_,
         action_reg_1__0_, action_reg_2__2_, action_reg_2__1_,
         action_reg_2__0_, action_reg_3__2_, action_reg_3__1_,
         action_reg_3__0_, action_reg_4__2_, action_reg_4__1_,
         action_reg_4__0_, action_reg_5__2_, action_reg_5__1_,
         action_reg_5__0_, action_reg_6__2_, action_reg_6__1_,
         action_reg_6__0_, action_reg_7__2_, action_reg_7__1_,
         action_reg_7__0_, in_valid_reg, N813, N814, start_write_flag, N1043,
         N1044, N1045, N1046, N1047, N1048, SRAM_192X32_WE,
         conv_sram_stop_flag_reg, SRAM_64X32_WE, N6115, N6116, N6117, N6118,
         N6119, N6120, N6121, N6122, N6123, N6124, N6125, N6126, N6127, N6128,
         N6129, N6130, N6291, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3404, n3405, n3415, n3416,
         mult_x_231_n48, mult_x_231_n39, mult_x_231_n11, mult_x_231_n10,
         mult_x_231_n9, mult_x_231_n8, mult_x_231_n7, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567,
         n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577,
         n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587,
         n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597,
         n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607,
         n3608, n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617,
         n3618, n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627,
         n3628, n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637,
         n3638, n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647,
         n3648, n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657,
         n3658, n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667,
         n3668, n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677,
         n3678, n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687,
         n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697,
         n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707,
         n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717,
         n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727,
         n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737,
         n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747,
         n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757,
         n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767,
         n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777,
         n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787,
         n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797,
         n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807,
         n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817,
         n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827,
         n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837,
         n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847,
         n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857,
         n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877,
         n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887,
         n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897,
         n3898, n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907,
         n3908, n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917,
         n3918, n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927,
         n3928, n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937,
         n3938, n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947,
         n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957,
         n3958, n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967,
         n3968, n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977,
         n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987,
         n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997,
         n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007,
         n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017,
         n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027,
         n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037,
         n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047,
         n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057,
         n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067,
         n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257,
         n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267,
         n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277,
         n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287,
         n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527,
         n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537,
         n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547,
         n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557,
         n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567,
         n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577,
         n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587,
         n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597,
         n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607,
         n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617,
         n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627,
         n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637,
         n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647,
         n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657,
         n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667,
         n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677,
         n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687,
         n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727,
         n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737,
         n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747,
         n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757,
         n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767,
         n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777,
         n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787,
         n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797,
         n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807,
         n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817,
         n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827,
         n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837,
         n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847,
         n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857,
         n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867,
         n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877,
         n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887,
         n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897,
         n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907,
         n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917,
         n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927,
         n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937,
         n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947,
         n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957,
         n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967,
         n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977,
         n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987,
         n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997,
         n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007,
         n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017,
         n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027,
         n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037,
         n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047,
         n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057,
         n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067,
         n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077,
         n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087,
         n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097,
         n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107,
         n6108, n6109, n6110, n6111, n6112, n6113, n6114, n61150, n61160,
         n61170, n61180, n61190, n61200, n61210, n61220, n61230, n61240,
         n61250, n61260, n61270, n61280, n61290, n61300, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n62910, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322;
  wire   [31:0] SRAM_192X32_out_decode;
  wire   [31:0] SRAM_64X32_in_decode;
  wire   [31:0] SRAM_64X32_out_decode;
  wire   [3:0] state;
  wire   [71:0] median_in;
  wire   [1:0] image_size_temp;
  wire   [8:0] cal_count;
  wire   [4:0] wait_conv_out_count;
  wire   [2:0] current_action_idx;
  wire   [3:0] action_idx;
  wire   [1:0] image_size_reg;
  wire   [7:0] SRAM_192X32_addr;
  wire   [2:0] set_count;
  wire   [3:0] template_count;
  wire   [71:0] template_reg;
  wire   [1:0] RGB_count;
  wire   [1:0] SRAM_192_32_in_count;
  wire   [7:0] max_temp;
  wire   [9:0] avg_temp;
  wire   [7:0] wgt_temp;
  wire   [31:0] gray_max_temp;
  wire   [31:0] gray_avg_reg;
  wire   [31:0] gray_wgt_reg;
  wire   [31:0] SRAM_192X32_data_in_reg;
  wire   [2:0] cal_count_5;
  wire   [7:6] rd_addr;
  wire   [7:0] wb_addr;
  wire   [31:0] SRAM_64X32_data_out;
  wire   [31:0] SRAM_192X32_data_out;
  wire   [3:0] cal_count_10;
  wire   [31:0] pool_temp;
  wire   [95:0] filter_result_reg;
  wire   [5:0] SRAM_64X32_addr;
  wire   [95:0] SRAM_out_buffer;
  wire   [7:0] median_result;
  wire   [15:0] product;
  wire   [19:0] conv_temp;
  wire   [19:0] conv_out_reg;
  wire   [2:0] conv_dly3;
  wire   [7:0] find_median_inst_final_mid;
  wire   [7:0] find_median_inst_min_pool_temp;
  wire   [7:0] find_median_inst_mid_mid_reg;
  wire   [7:0] find_median_inst_max_min_reg;
  wire   [7:0] find_median_inst_min_max;
  wire   [7:0] find_median_inst_min3_reg;
  wire   [7:0] find_median_inst_min2_reg;
  wire   [7:0] find_median_inst_min1_reg;
  wire   [7:0] find_median_inst_mid_mid;
  wire   [7:0] find_median_inst_mid3_reg;
  wire   [7:0] find_median_inst_mid2_reg;
  wire   [7:0] find_median_inst_mid1_reg;
  wire   [7:0] find_median_inst_max_min;
  wire   [7:0] find_median_inst_max3_reg;
  wire   [7:0] find_median_inst_max2_reg;
  wire   [7:0] find_median_inst_max1_reg;
  wire   [7:0] find_median_inst_max3;
  wire   [7:0] find_median_inst_mid3;
  wire   [7:0] find_median_inst_min3;
  wire   [7:0] find_median_inst_max2;
  wire   [7:0] find_median_inst_mid2;
  wire   [7:0] find_median_inst_min2;
  wire   [7:0] find_median_inst_max1;
  wire   [7:0] find_median_inst_mid1;
  wire   [7:0] find_median_inst_min1;

  SRAM_192X32 SRAM_192_32_inst_SRAM_192X32_inst ( .A0(SRAM_192X32_addr[0]), 
        .A1(SRAM_192X32_addr[1]), .A2(SRAM_192X32_addr[2]), .A3(
        SRAM_192X32_addr[3]), .A4(SRAM_192X32_addr[4]), .A5(
        SRAM_192X32_addr[5]), .A6(SRAM_192X32_addr[6]), .A7(
        SRAM_192X32_addr[7]), .CK(clk), .CS(n2863), .DI0(
        SRAM_192X32_data_in_reg[0]), .DI1(SRAM_192X32_data_in_reg[1]), .DI10(
        SRAM_192X32_data_in_reg[10]), .DI11(SRAM_192X32_data_in_reg[11]), 
        .DI12(SRAM_192X32_data_in_reg[12]), .DI13(SRAM_192X32_data_in_reg[13]), 
        .DI14(SRAM_192X32_data_in_reg[14]), .DI15(SRAM_192X32_data_in_reg[15]), 
        .DI16(SRAM_192X32_data_in_reg[16]), .DI17(SRAM_192X32_data_in_reg[17]), 
        .DI18(SRAM_192X32_data_in_reg[18]), .DI19(SRAM_192X32_data_in_reg[19]), 
        .DI2(SRAM_192X32_data_in_reg[2]), .DI20(SRAM_192X32_data_in_reg[20]), 
        .DI21(SRAM_192X32_data_in_reg[21]), .DI22(SRAM_192X32_data_in_reg[22]), 
        .DI23(SRAM_192X32_data_in_reg[23]), .DI24(SRAM_192X32_data_in_reg[24]), 
        .DI25(SRAM_192X32_data_in_reg[25]), .DI26(SRAM_192X32_data_in_reg[26]), 
        .DI27(SRAM_192X32_data_in_reg[27]), .DI28(SRAM_192X32_data_in_reg[28]), 
        .DI29(SRAM_192X32_data_in_reg[29]), .DI3(SRAM_192X32_data_in_reg[3]), 
        .DI30(SRAM_192X32_data_in_reg[30]), .DI31(SRAM_192X32_data_in_reg[31]), 
        .DI4(SRAM_192X32_data_in_reg[4]), .DI5(SRAM_192X32_data_in_reg[5]), 
        .DI6(SRAM_192X32_data_in_reg[6]), .DI7(SRAM_192X32_data_in_reg[7]), 
        .DI8(SRAM_192X32_data_in_reg[8]), .DI9(SRAM_192X32_data_in_reg[9]), 
        .OE(n2863), .WEB(n3415), .DO0(SRAM_192X32_data_out[0]), .DO1(
        SRAM_192X32_data_out[1]), .DO10(SRAM_192X32_data_out[10]), .DO11(
        SRAM_192X32_data_out[11]), .DO12(SRAM_192X32_data_out[12]), .DO13(
        SRAM_192X32_data_out[13]), .DO14(SRAM_192X32_data_out[14]), .DO15(
        SRAM_192X32_data_out[15]), .DO16(SRAM_192X32_data_out[16]), .DO17(
        SRAM_192X32_data_out[17]), .DO18(SRAM_192X32_data_out[18]), .DO19(
        SRAM_192X32_data_out[19]), .DO2(SRAM_192X32_data_out[2]), .DO20(
        SRAM_192X32_data_out[20]), .DO21(SRAM_192X32_data_out[21]), .DO22(
        SRAM_192X32_data_out[22]), .DO23(SRAM_192X32_data_out[23]), .DO24(
        SRAM_192X32_data_out[24]), .DO25(SRAM_192X32_data_out[25]), .DO26(
        SRAM_192X32_data_out[26]), .DO27(SRAM_192X32_data_out[27]), .DO28(
        SRAM_192X32_data_out[28]), .DO29(SRAM_192X32_data_out[29]), .DO3(
        SRAM_192X32_data_out[3]), .DO30(SRAM_192X32_data_out[30]), .DO31(
        SRAM_192X32_data_out[31]), .DO4(SRAM_192X32_data_out[4]), .DO5(
        SRAM_192X32_data_out[5]), .DO6(SRAM_192X32_data_out[6]), .DO7(
        SRAM_192X32_data_out[7]), .DO8(SRAM_192X32_data_out[8]), .DO9(
        SRAM_192X32_data_out[9]) );
  SRAM_64X32 SRAM_64_32_inst_SRAM_64X32_inst ( .A0(SRAM_64X32_addr[0]), .A1(
        SRAM_64X32_addr[1]), .A2(SRAM_64X32_addr[2]), .A3(SRAM_64X32_addr[3]), 
        .A4(SRAM_64X32_addr[4]), .A5(SRAM_64X32_addr[5]), .CK(clk), .CS(n2863), 
        .DI0(SRAM_64X32_in_decode[0]), .DI1(SRAM_64X32_in_decode[1]), .DI10(
        SRAM_64X32_in_decode[10]), .DI11(SRAM_64X32_in_decode[11]), .DI12(
        SRAM_64X32_in_decode[12]), .DI13(SRAM_64X32_in_decode[13]), .DI14(
        SRAM_64X32_in_decode[14]), .DI15(SRAM_64X32_in_decode[15]), .DI16(
        SRAM_64X32_in_decode[16]), .DI17(SRAM_64X32_in_decode[17]), .DI18(
        SRAM_64X32_in_decode[18]), .DI19(SRAM_64X32_in_decode[19]), .DI2(
        SRAM_64X32_in_decode[2]), .DI20(SRAM_64X32_in_decode[20]), .DI21(
        SRAM_64X32_in_decode[21]), .DI22(SRAM_64X32_in_decode[22]), .DI23(
        SRAM_64X32_in_decode[23]), .DI24(SRAM_64X32_in_decode[24]), .DI25(
        SRAM_64X32_in_decode[25]), .DI26(SRAM_64X32_in_decode[26]), .DI27(
        SRAM_64X32_in_decode[27]), .DI28(SRAM_64X32_in_decode[28]), .DI29(
        SRAM_64X32_in_decode[29]), .DI3(SRAM_64X32_in_decode[3]), .DI30(
        SRAM_64X32_in_decode[30]), .DI31(SRAM_64X32_in_decode[31]), .DI4(
        SRAM_64X32_in_decode[4]), .DI5(SRAM_64X32_in_decode[5]), .DI6(
        SRAM_64X32_in_decode[6]), .DI7(SRAM_64X32_in_decode[7]), .DI8(
        SRAM_64X32_in_decode[8]), .DI9(SRAM_64X32_in_decode[9]), .OE(n2863), 
        .WEB(n3416), .DO0(SRAM_64X32_data_out[0]), .DO1(SRAM_64X32_data_out[1]), .DO10(SRAM_64X32_data_out[10]), .DO11(SRAM_64X32_data_out[11]), .DO12(
        SRAM_64X32_data_out[12]), .DO13(SRAM_64X32_data_out[13]), .DO14(
        SRAM_64X32_data_out[14]), .DO15(SRAM_64X32_data_out[15]), .DO16(
        SRAM_64X32_data_out[16]), .DO17(SRAM_64X32_data_out[17]), .DO18(
        SRAM_64X32_data_out[18]), .DO19(SRAM_64X32_data_out[19]), .DO2(
        SRAM_64X32_data_out[2]), .DO20(SRAM_64X32_data_out[20]), .DO21(
        SRAM_64X32_data_out[21]), .DO22(SRAM_64X32_data_out[22]), .DO23(
        SRAM_64X32_data_out[23]), .DO24(SRAM_64X32_data_out[24]), .DO25(
        SRAM_64X32_data_out[25]), .DO26(SRAM_64X32_data_out[26]), .DO27(
        SRAM_64X32_data_out[27]), .DO28(SRAM_64X32_data_out[28]), .DO29(
        SRAM_64X32_data_out[29]), .DO3(SRAM_64X32_data_out[3]), .DO30(
        SRAM_64X32_data_out[30]), .DO31(SRAM_64X32_data_out[31]), .DO4(
        SRAM_64X32_data_out[4]), .DO5(SRAM_64X32_data_out[5]), .DO6(
        SRAM_64X32_data_out[6]), .DO7(SRAM_64X32_data_out[7]), .DO8(
        SRAM_64X32_data_out[8]), .DO9(SRAM_64X32_data_out[9]) );
  QDFFS in_valid_reg_reg ( .D(n3493), .CK(clk), .Q(in_valid_reg) );
  QDFFS template_reg_reg_7__0_ ( .D(n3334), .CK(clk), .Q(template_reg[8]) );
  QDFFS template_reg_reg_7__7_ ( .D(n3333), .CK(clk), .Q(template_reg[15]) );
  QDFFS template_reg_reg_7__6_ ( .D(n3332), .CK(clk), .Q(template_reg[14]) );
  QDFFS template_reg_reg_7__5_ ( .D(n3331), .CK(clk), .Q(template_reg[13]) );
  QDFFS template_reg_reg_7__4_ ( .D(n3330), .CK(clk), .Q(template_reg[12]) );
  QDFFS template_reg_reg_7__3_ ( .D(n3329), .CK(clk), .Q(template_reg[11]) );
  QDFFS template_reg_reg_7__2_ ( .D(n3328), .CK(clk), .Q(template_reg[10]) );
  QDFFS template_reg_reg_7__1_ ( .D(n3327), .CK(clk), .Q(template_reg[9]) );
  QDFFS template_reg_reg_3__0_ ( .D(n3302), .CK(clk), .Q(template_reg[40]) );
  QDFFS template_reg_reg_3__7_ ( .D(n3301), .CK(clk), .Q(template_reg[47]) );
  QDFFS template_reg_reg_3__6_ ( .D(n3300), .CK(clk), .Q(template_reg[46]) );
  QDFFS template_reg_reg_3__5_ ( .D(n3299), .CK(clk), .Q(template_reg[45]) );
  QDFFS template_reg_reg_3__4_ ( .D(n3298), .CK(clk), .Q(template_reg[44]) );
  QDFFS template_reg_reg_3__3_ ( .D(n3297), .CK(clk), .Q(template_reg[43]) );
  QDFFS template_reg_reg_3__2_ ( .D(n3296), .CK(clk), .Q(template_reg[42]) );
  QDFFS template_reg_reg_3__1_ ( .D(n3295), .CK(clk), .Q(template_reg[41]) );
  QDFFS template_reg_reg_5__0_ ( .D(n3318), .CK(clk), .Q(template_reg[24]) );
  QDFFS template_reg_reg_5__7_ ( .D(n3317), .CK(clk), .Q(template_reg[31]) );
  QDFFS template_reg_reg_5__6_ ( .D(n3316), .CK(clk), .Q(template_reg[30]) );
  QDFFS template_reg_reg_5__5_ ( .D(n3315), .CK(clk), .Q(template_reg[29]) );
  QDFFS template_reg_reg_5__4_ ( .D(n3314), .CK(clk), .Q(template_reg[28]) );
  QDFFS template_reg_reg_5__3_ ( .D(n3313), .CK(clk), .Q(template_reg[27]) );
  QDFFS template_reg_reg_5__2_ ( .D(n3312), .CK(clk), .Q(template_reg[26]) );
  QDFFS template_reg_reg_5__1_ ( .D(n3311), .CK(clk), .Q(template_reg[25]) );
  QDFFS template_reg_reg_1__0_ ( .D(n3286), .CK(clk), .Q(template_reg[56]) );
  QDFFS template_reg_reg_1__7_ ( .D(n3285), .CK(clk), .Q(template_reg[63]) );
  QDFFS template_reg_reg_1__6_ ( .D(n3284), .CK(clk), .Q(template_reg[62]) );
  QDFFS template_reg_reg_1__5_ ( .D(n3283), .CK(clk), .Q(template_reg[61]) );
  QDFFS template_reg_reg_1__4_ ( .D(n3282), .CK(clk), .Q(template_reg[60]) );
  QDFFS template_reg_reg_1__3_ ( .D(n3281), .CK(clk), .Q(template_reg[59]) );
  QDFFS template_reg_reg_1__2_ ( .D(n3280), .CK(clk), .Q(template_reg[58]) );
  QDFFS template_reg_reg_1__1_ ( .D(n3279), .CK(clk), .Q(template_reg[57]) );
  QDFFS template_reg_reg_6__0_ ( .D(n3326), .CK(clk), .Q(template_reg[16]) );
  QDFFS template_reg_reg_6__7_ ( .D(n3325), .CK(clk), .Q(template_reg[23]) );
  QDFFS template_reg_reg_6__6_ ( .D(n3324), .CK(clk), .Q(template_reg[22]) );
  QDFFS template_reg_reg_6__5_ ( .D(n3323), .CK(clk), .Q(template_reg[21]) );
  QDFFS template_reg_reg_6__4_ ( .D(n3322), .CK(clk), .Q(template_reg[20]) );
  QDFFS template_reg_reg_6__3_ ( .D(n3321), .CK(clk), .Q(template_reg[19]) );
  QDFFS template_reg_reg_6__2_ ( .D(n3320), .CK(clk), .Q(template_reg[18]) );
  QDFFS template_reg_reg_6__1_ ( .D(n3319), .CK(clk), .Q(template_reg[17]) );
  QDFFS template_reg_reg_4__0_ ( .D(n3310), .CK(clk), .Q(template_reg[32]) );
  QDFFS template_reg_reg_4__7_ ( .D(n3309), .CK(clk), .Q(template_reg[39]) );
  QDFFS template_reg_reg_4__6_ ( .D(n3308), .CK(clk), .Q(template_reg[38]) );
  QDFFS template_reg_reg_4__5_ ( .D(n3307), .CK(clk), .Q(template_reg[37]) );
  QDFFS template_reg_reg_4__4_ ( .D(n3306), .CK(clk), .Q(template_reg[36]) );
  QDFFS template_reg_reg_4__3_ ( .D(n3305), .CK(clk), .Q(template_reg[35]) );
  QDFFS template_reg_reg_4__2_ ( .D(n3304), .CK(clk), .Q(template_reg[34]) );
  QDFFS template_reg_reg_4__1_ ( .D(n3303), .CK(clk), .Q(template_reg[33]) );
  QDFFS template_reg_reg_2__0_ ( .D(n3294), .CK(clk), .Q(template_reg[48]) );
  QDFFS template_reg_reg_2__7_ ( .D(n3293), .CK(clk), .Q(template_reg[55]) );
  QDFFS template_reg_reg_2__6_ ( .D(n3292), .CK(clk), .Q(template_reg[54]) );
  QDFFS template_reg_reg_2__5_ ( .D(n3291), .CK(clk), .Q(template_reg[53]) );
  QDFFS template_reg_reg_2__4_ ( .D(n3290), .CK(clk), .Q(template_reg[52]) );
  QDFFS template_reg_reg_2__3_ ( .D(n3289), .CK(clk), .Q(template_reg[51]) );
  QDFFS template_reg_reg_2__2_ ( .D(n3288), .CK(clk), .Q(template_reg[50]) );
  QDFFS template_reg_reg_2__1_ ( .D(n3287), .CK(clk), .Q(template_reg[49]) );
  QDFFS template_reg_reg_8__0_ ( .D(n3342), .CK(clk), .Q(template_reg[0]) );
  QDFFS template_reg_reg_8__7_ ( .D(n3341), .CK(clk), .Q(template_reg[7]) );
  QDFFS template_reg_reg_8__6_ ( .D(n3340), .CK(clk), .Q(template_reg[6]) );
  QDFFS template_reg_reg_8__5_ ( .D(n3339), .CK(clk), .Q(template_reg[5]) );
  QDFFS template_reg_reg_8__4_ ( .D(n3338), .CK(clk), .Q(template_reg[4]) );
  QDFFS template_reg_reg_8__3_ ( .D(n3337), .CK(clk), .Q(template_reg[3]) );
  QDFFS template_reg_reg_8__2_ ( .D(n3336), .CK(clk), .Q(template_reg[2]) );
  QDFFS template_reg_reg_8__1_ ( .D(n3335), .CK(clk), .Q(template_reg[1]) );
  QDFFS template_reg_reg_0__0_ ( .D(n3278), .CK(clk), .Q(template_reg[64]) );
  QDFFS template_reg_reg_0__7_ ( .D(n3277), .CK(clk), .Q(template_reg[71]) );
  QDFFS template_reg_reg_0__6_ ( .D(n3276), .CK(clk), .Q(template_reg[70]) );
  QDFFS template_reg_reg_0__5_ ( .D(n3275), .CK(clk), .Q(template_reg[69]) );
  QDFFS template_reg_reg_0__4_ ( .D(n3274), .CK(clk), .Q(template_reg[68]) );
  QDFFS template_reg_reg_0__3_ ( .D(n3273), .CK(clk), .Q(template_reg[67]) );
  QDFFS template_reg_reg_0__2_ ( .D(n3272), .CK(clk), .Q(template_reg[66]) );
  QDFFS template_reg_reg_0__1_ ( .D(n3271), .CK(clk), .Q(template_reg[65]) );
  QDFFS product_reg_14_ ( .D(N6129), .CK(clk), .Q(product[14]) );
  QDFFS product_reg_13_ ( .D(N6128), .CK(clk), .Q(product[13]) );
  QDFFS product_reg_12_ ( .D(N6127), .CK(clk), .Q(product[12]) );
  QDFFS product_reg_11_ ( .D(N6126), .CK(clk), .Q(product[11]) );
  QDFFS product_reg_10_ ( .D(N6125), .CK(clk), .Q(product[10]) );
  QDFFS product_reg_9_ ( .D(N6124), .CK(clk), .Q(product[9]) );
  QDFFS product_reg_8_ ( .D(N6123), .CK(clk), .Q(product[8]) );
  QDFFS product_reg_7_ ( .D(N6122), .CK(clk), .Q(product[7]) );
  QDFFS product_reg_6_ ( .D(N6121), .CK(clk), .Q(product[6]) );
  QDFFS product_reg_5_ ( .D(N6120), .CK(clk), .Q(product[5]) );
  QDFFS product_reg_4_ ( .D(N6119), .CK(clk), .Q(product[4]) );
  QDFFS product_reg_3_ ( .D(N6118), .CK(clk), .Q(product[3]) );
  QDFFS product_reg_2_ ( .D(N6117), .CK(clk), .Q(product[2]) );
  QDFFS product_reg_1_ ( .D(N6116), .CK(clk), .Q(product[1]) );
  QDFFS product_reg_0_ ( .D(N6115), .CK(clk), .Q(product[0]) );
  QDFFS action_reg_reg_6__0_ ( .D(n3391), .CK(clk), .Q(action_reg_6__0_) );
  QDFFS action_reg_reg_6__2_ ( .D(n3390), .CK(clk), .Q(action_reg_6__2_) );
  QDFFS action_reg_reg_6__1_ ( .D(n3389), .CK(clk), .Q(action_reg_6__1_) );
  QDFFS action_reg_reg_4__0_ ( .D(n3385), .CK(clk), .Q(action_reg_4__0_) );
  QDFFS action_reg_reg_4__2_ ( .D(n3384), .CK(clk), .Q(action_reg_4__2_) );
  QDFFS action_reg_reg_4__1_ ( .D(n3383), .CK(clk), .Q(action_reg_4__1_) );
  QDFFS action_reg_reg_7__0_ ( .D(n3394), .CK(clk), .Q(action_reg_7__0_) );
  QDFFS action_reg_reg_7__2_ ( .D(n3393), .CK(clk), .Q(action_reg_7__2_) );
  QDFFS action_reg_reg_7__1_ ( .D(n3392), .CK(clk), .Q(action_reg_7__1_) );
  QDFFS action_reg_reg_5__0_ ( .D(n3388), .CK(clk), .Q(action_reg_5__0_) );
  QDFFS action_reg_reg_5__2_ ( .D(n3387), .CK(clk), .Q(action_reg_5__2_) );
  QDFFS action_reg_reg_5__1_ ( .D(n3386), .CK(clk), .Q(action_reg_5__1_) );
  QDFFS action_reg_reg_3__0_ ( .D(n3382), .CK(clk), .Q(action_reg_3__0_) );
  QDFFS action_reg_reg_3__2_ ( .D(n3381), .CK(clk), .Q(action_reg_3__2_) );
  QDFFS action_reg_reg_3__1_ ( .D(n3380), .CK(clk), .Q(action_reg_3__1_) );
  QDFFS action_reg_reg_1__0_ ( .D(n3376), .CK(clk), .Q(action_reg_1__0_) );
  QDFFS action_reg_reg_1__2_ ( .D(n3375), .CK(clk), .Q(action_reg_1__2_) );
  QDFFS action_reg_reg_1__1_ ( .D(n3374), .CK(clk), .Q(action_reg_1__1_) );
  QDFFS action_reg_reg_0__0_ ( .D(n3373), .CK(clk), .Q(action_reg_0__0_) );
  QDFFS action_reg_reg_0__1_ ( .D(n3372), .CK(clk), .Q(action_reg_0__1_) );
  QDFFS action_reg_reg_2__0_ ( .D(n3379), .CK(clk), .Q(action_reg_2__0_) );
  QDFFS action_reg_reg_2__2_ ( .D(n3378), .CK(clk), .Q(action_reg_2__2_) );
  QDFFS action_reg_reg_2__1_ ( .D(n3377), .CK(clk), .Q(action_reg_2__1_) );
  QDFFS SRAM_192X32_data_in_reg_reg_0_ ( .D(n3267), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[0]) );
  QDFFS SRAM_192X32_data_in_reg_reg_1_ ( .D(n3266), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[1]) );
  QDFFS SRAM_192X32_data_in_reg_reg_2_ ( .D(n3265), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[2]) );
  QDFFS SRAM_192X32_data_in_reg_reg_3_ ( .D(n3264), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[3]) );
  QDFFS SRAM_192X32_data_in_reg_reg_4_ ( .D(n3263), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[4]) );
  QDFFS SRAM_192X32_data_in_reg_reg_5_ ( .D(n3262), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[5]) );
  QDFFS SRAM_192X32_data_in_reg_reg_6_ ( .D(n3261), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[6]) );
  QDFFS SRAM_192X32_data_in_reg_reg_7_ ( .D(n3260), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[7]) );
  QDFFS SRAM_192X32_data_in_reg_reg_8_ ( .D(n3259), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[8]) );
  QDFFS SRAM_192X32_data_in_reg_reg_9_ ( .D(n3258), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[9]) );
  QDFFS SRAM_192X32_data_in_reg_reg_10_ ( .D(n3257), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[10]) );
  QDFFS SRAM_192X32_data_in_reg_reg_11_ ( .D(n3256), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[11]) );
  QDFFS SRAM_192X32_data_in_reg_reg_12_ ( .D(n3255), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[12]) );
  QDFFS SRAM_192X32_data_in_reg_reg_13_ ( .D(n3254), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[13]) );
  QDFFS SRAM_192X32_data_in_reg_reg_14_ ( .D(n3253), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[14]) );
  QDFFS SRAM_192X32_data_in_reg_reg_15_ ( .D(n3252), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[15]) );
  QDFFS SRAM_192X32_data_in_reg_reg_16_ ( .D(n3251), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[16]) );
  QDFFS SRAM_192X32_data_in_reg_reg_17_ ( .D(n3250), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[17]) );
  QDFFS SRAM_192X32_data_in_reg_reg_18_ ( .D(n3249), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[18]) );
  QDFFS SRAM_192X32_data_in_reg_reg_19_ ( .D(n3248), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[19]) );
  QDFFS SRAM_192X32_data_in_reg_reg_20_ ( .D(n3247), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[20]) );
  QDFFS SRAM_192X32_data_in_reg_reg_21_ ( .D(n3246), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[21]) );
  QDFFS SRAM_192X32_data_in_reg_reg_22_ ( .D(n3245), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[22]) );
  QDFFS SRAM_192X32_data_in_reg_reg_23_ ( .D(n3244), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[23]) );
  QDFFS SRAM_192X32_data_in_reg_reg_24_ ( .D(n3243), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[24]) );
  QDFFS SRAM_192X32_data_in_reg_reg_25_ ( .D(n3242), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[25]) );
  QDFFS SRAM_192X32_data_in_reg_reg_26_ ( .D(n3241), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[26]) );
  QDFFS SRAM_192X32_data_in_reg_reg_27_ ( .D(n3240), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[27]) );
  QDFFS SRAM_192X32_data_in_reg_reg_28_ ( .D(n3239), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[28]) );
  QDFFS SRAM_192X32_data_in_reg_reg_29_ ( .D(n3238), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[29]) );
  QDFFS SRAM_192X32_data_in_reg_reg_30_ ( .D(n3237), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[30]) );
  QDFFS SRAM_192X32_data_in_reg_reg_31_ ( .D(n3236), .CK(clk), .Q(
        SRAM_192X32_data_in_reg[31]) );
  QDFFS filter_result_reg_reg_0__3__7_ ( .D(n3167), .CK(clk), .Q(
        filter_result_reg[71]) );
  QDFFS filter_result_reg_reg_0__2__7_ ( .D(n3166), .CK(clk), .Q(
        filter_result_reg[79]) );
  QDFFS filter_result_reg_reg_0__1__7_ ( .D(n3165), .CK(clk), .Q(
        filter_result_reg[87]) );
  QDFFS filter_result_reg_reg_0__0__7_ ( .D(n3164), .CK(clk), .Q(
        filter_result_reg[95]) );
  QDFFS SRAM_64X32_data_in_reg_reg_31_ ( .D(n3163), .CK(clk), .Q(
        SRAM_64X32_in_decode[31]) );
  QDFFS SRAM_out_buffer_reg_1__3__7_ ( .D(n3141), .CK(clk), .Q(
        SRAM_out_buffer[39]) );
  QDFFS SRAM_out_buffer_reg_0__3__7_ ( .D(n3140), .CK(clk), .Q(
        SRAM_out_buffer[71]) );
  QDFFS SRAM_out_buffer_reg_2__3__7_ ( .D(n3139), .CK(clk), .Q(
        SRAM_out_buffer[7]) );
  QDFFS SRAM_out_buffer_reg_1__0__7_ ( .D(n2926), .CK(clk), .Q(
        SRAM_out_buffer[63]) );
  QDFFS SRAM_out_buffer_reg_0__0__7_ ( .D(n2925), .CK(clk), .Q(
        SRAM_out_buffer[95]) );
  QDFFS SRAM_out_buffer_reg_2__0__7_ ( .D(n2887), .CK(clk), .Q(
        SRAM_out_buffer[31]) );
  QDFFS SRAM_out_buffer_reg_1__3__6_ ( .D(n3144), .CK(clk), .Q(
        SRAM_out_buffer[38]) );
  QDFFS SRAM_out_buffer_reg_0__3__6_ ( .D(n3143), .CK(clk), .Q(
        SRAM_out_buffer[70]) );
  QDFFS SRAM_out_buffer_reg_2__3__6_ ( .D(n3142), .CK(clk), .Q(
        SRAM_out_buffer[6]) );
  QDFFS SRAM_out_buffer_reg_1__0__6_ ( .D(n2938), .CK(clk), .Q(
        SRAM_out_buffer[62]) );
  QDFFS SRAM_out_buffer_reg_0__0__6_ ( .D(n2937), .CK(clk), .Q(
        SRAM_out_buffer[94]) );
  QDFFS SRAM_out_buffer_reg_2__0__6_ ( .D(n2930), .CK(clk), .Q(
        SRAM_out_buffer[30]) );
  QDFFS SRAM_out_buffer_reg_1__3__5_ ( .D(n3147), .CK(clk), .Q(
        SRAM_out_buffer[37]) );
  QDFFS SRAM_out_buffer_reg_0__3__5_ ( .D(n3146), .CK(clk), .Q(
        SRAM_out_buffer[69]) );
  QDFFS SRAM_out_buffer_reg_2__3__5_ ( .D(n3145), .CK(clk), .Q(
        SRAM_out_buffer[5]) );
  QDFFS SRAM_out_buffer_reg_1__0__5_ ( .D(n2950), .CK(clk), .Q(
        SRAM_out_buffer[61]) );
  QDFFS SRAM_out_buffer_reg_0__0__5_ ( .D(n2949), .CK(clk), .Q(
        SRAM_out_buffer[93]) );
  QDFFS SRAM_out_buffer_reg_2__0__5_ ( .D(n2942), .CK(clk), .Q(
        SRAM_out_buffer[29]) );
  QDFFS SRAM_out_buffer_reg_1__3__4_ ( .D(n3150), .CK(clk), .Q(
        SRAM_out_buffer[36]) );
  QDFFS SRAM_out_buffer_reg_0__3__4_ ( .D(n3149), .CK(clk), .Q(
        SRAM_out_buffer[68]) );
  QDFFS SRAM_out_buffer_reg_2__3__4_ ( .D(n3148), .CK(clk), .Q(
        SRAM_out_buffer[4]) );
  QDFFS SRAM_out_buffer_reg_1__0__4_ ( .D(n2962), .CK(clk), .Q(
        SRAM_out_buffer[60]) );
  QDFFS SRAM_out_buffer_reg_0__0__4_ ( .D(n2961), .CK(clk), .Q(
        SRAM_out_buffer[92]) );
  QDFFS SRAM_out_buffer_reg_2__0__4_ ( .D(n2954), .CK(clk), .Q(
        SRAM_out_buffer[28]) );
  QDFFS SRAM_out_buffer_reg_1__3__3_ ( .D(n3153), .CK(clk), .Q(
        SRAM_out_buffer[35]) );
  QDFFS SRAM_out_buffer_reg_0__3__3_ ( .D(n3152), .CK(clk), .Q(
        SRAM_out_buffer[67]) );
  QDFFS SRAM_out_buffer_reg_2__3__3_ ( .D(n3151), .CK(clk), .Q(
        SRAM_out_buffer[3]) );
  QDFFS SRAM_out_buffer_reg_1__0__3_ ( .D(n2974), .CK(clk), .Q(
        SRAM_out_buffer[59]) );
  QDFFS SRAM_out_buffer_reg_0__0__3_ ( .D(n2973), .CK(clk), .Q(
        SRAM_out_buffer[91]) );
  QDFFS SRAM_out_buffer_reg_2__0__3_ ( .D(n2966), .CK(clk), .Q(
        SRAM_out_buffer[27]) );
  QDFFS SRAM_out_buffer_reg_1__3__2_ ( .D(n3156), .CK(clk), .Q(
        SRAM_out_buffer[34]) );
  QDFFS SRAM_out_buffer_reg_0__3__2_ ( .D(n3155), .CK(clk), .Q(
        SRAM_out_buffer[66]) );
  QDFFS SRAM_out_buffer_reg_2__3__2_ ( .D(n3154), .CK(clk), .Q(
        SRAM_out_buffer[2]) );
  QDFFS SRAM_out_buffer_reg_1__0__2_ ( .D(n2986), .CK(clk), .Q(
        SRAM_out_buffer[58]) );
  QDFFS SRAM_out_buffer_reg_0__0__2_ ( .D(n2985), .CK(clk), .Q(
        SRAM_out_buffer[90]) );
  QDFFS SRAM_out_buffer_reg_2__0__2_ ( .D(n2978), .CK(clk), .Q(
        SRAM_out_buffer[26]) );
  QDFFS SRAM_out_buffer_reg_1__2__1_ ( .D(n3132), .CK(clk), .Q(
        SRAM_out_buffer[41]) );
  QDFFS SRAM_out_buffer_reg_0__2__1_ ( .D(n3131), .CK(clk), .Q(
        SRAM_out_buffer[73]) );
  QDFFS SRAM_out_buffer_reg_2__2__1_ ( .D(n3128), .CK(clk), .Q(
        SRAM_out_buffer[9]) );
  QDFFS SRAM_out_buffer_reg_1__1__1_ ( .D(n3052), .CK(clk), .Q(
        SRAM_out_buffer[49]) );
  QDFFS SRAM_out_buffer_reg_0__1__1_ ( .D(n3051), .CK(clk), .Q(
        SRAM_out_buffer[81]) );
  QDFFS SRAM_out_buffer_reg_2__1__1_ ( .D(n3048), .CK(clk), .Q(
        SRAM_out_buffer[17]) );
  QDFFS SRAM_out_buffer_reg_1__2__0_ ( .D(n3138), .CK(clk), .Q(
        SRAM_out_buffer[40]) );
  QDFFS SRAM_out_buffer_reg_0__2__0_ ( .D(n3137), .CK(clk), .Q(
        SRAM_out_buffer[72]) );
  QDFFS SRAM_out_buffer_reg_2__2__0_ ( .D(n3134), .CK(clk), .Q(
        SRAM_out_buffer[8]) );
  QDFFS SRAM_out_buffer_reg_1__1__0_ ( .D(n3058), .CK(clk), .Q(
        SRAM_out_buffer[48]) );
  QDFFS SRAM_out_buffer_reg_0__1__0_ ( .D(n3057), .CK(clk), .Q(
        SRAM_out_buffer[80]) );
  QDFFS SRAM_out_buffer_reg_2__1__0_ ( .D(n3054), .CK(clk), .Q(
        SRAM_out_buffer[16]) );
  QDFFS SRAM_out_buffer_reg_1__2__7_ ( .D(n3096), .CK(clk), .Q(
        SRAM_out_buffer[47]) );
  QDFFS SRAM_out_buffer_reg_0__2__7_ ( .D(n3095), .CK(clk), .Q(
        SRAM_out_buffer[79]) );
  QDFFS window_reg_1__4__7_ ( .D(n3094), .CK(clk), .Q(window_1__4__7_) );
  QDFFS window_reg_0__4__7_ ( .D(n3093), .CK(clk), .Q(window_0__4__7_) );
  QDFFS pool_temp_reg_1__7_ ( .D(n3092), .CK(clk), .Q(pool_temp[23]) );
  QDFFS SRAM_64X32_data_in_reg_reg_23_ ( .D(n3091), .CK(clk), .Q(
        SRAM_64X32_in_decode[23]) );
  QDFFS pool_temp_reg_3__7_ ( .D(n3076), .CK(clk), .Q(pool_temp[7]) );
  QDFFS SRAM_64X32_data_in_reg_reg_7_ ( .D(n3075), .CK(clk), .Q(
        SRAM_64X32_in_decode[7]) );
  QDFFS SRAM_out_buffer_reg_2__2__7_ ( .D(n3060), .CK(clk), .Q(
        SRAM_out_buffer[15]) );
  QDFFS window_reg_2__4__7_ ( .D(n3059), .CK(clk), .Q(window_2__4__7_) );
  QDFFS SRAM_out_buffer_reg_1__1__7_ ( .D(n3016), .CK(clk), .Q(
        SRAM_out_buffer[55]) );
  QDFFS SRAM_out_buffer_reg_0__1__7_ ( .D(n3015), .CK(clk), .Q(
        SRAM_out_buffer[87]) );
  QDFFS window_reg_1__3__7_ ( .D(n3014), .CK(clk), .Q(window_1__3__7_) );
  QDFFS window_reg_0__3__7_ ( .D(n3013), .CK(clk), .Q(window_0__3__7_) );
  QDFFS window_reg_1__2__7_ ( .D(n2924), .CK(clk), .Q(median_in[31]) );
  QDFFS window_reg_1__1__7_ ( .D(n2923), .CK(clk), .Q(median_in[39]) );
  QDFFS window_reg_1__0__7_ ( .D(n2922), .CK(clk), .Q(median_in[47]) );
  QDFFS window_reg_0__2__7_ ( .D(n2921), .CK(clk), .Q(median_in[55]) );
  QDFFS window_reg_0__1__7_ ( .D(n2920), .CK(clk), .Q(median_in[63]) );
  QDFFS window_reg_0__0__7_ ( .D(n2919), .CK(clk), .Q(median_in[71]) );
  QDFFS SRAM_out_buffer_reg_2__1__7_ ( .D(n3012), .CK(clk), .Q(
        SRAM_out_buffer[23]) );
  QDFFS window_reg_2__3__7_ ( .D(n3011), .CK(clk), .Q(window_2__3__7_) );
  QDFFS pool_temp_reg_0__7_ ( .D(n2918), .CK(clk), .Q(pool_temp[31]) );
  QDFFS pool_temp_reg_2__7_ ( .D(n2903), .CK(clk), .Q(pool_temp[15]) );
  QDFFS SRAM_64X32_data_in_reg_reg_15_ ( .D(n2902), .CK(clk), .Q(
        SRAM_64X32_in_decode[15]) );
  QDFFS window_reg_2__2__7_ ( .D(n2886), .CK(clk), .Q(median_in[7]) );
  QDFFS window_reg_2__1__7_ ( .D(n2885), .CK(clk), .Q(median_in[15]) );
  QDFFS window_reg_2__0__7_ ( .D(n2884), .CK(clk), .Q(median_in[23]) );
  QDFFS SRAM_out_buffer_reg_1__2__6_ ( .D(n3102), .CK(clk), .Q(
        SRAM_out_buffer[46]) );
  QDFFS SRAM_out_buffer_reg_0__2__6_ ( .D(n3101), .CK(clk), .Q(
        SRAM_out_buffer[78]) );
  QDFFS window_reg_1__4__6_ ( .D(n3100), .CK(clk), .Q(window_1__4__6_) );
  QDFFS window_reg_0__4__6_ ( .D(n3099), .CK(clk), .Q(window_0__4__6_) );
  QDFFS SRAM_out_buffer_reg_2__2__6_ ( .D(n3098), .CK(clk), .Q(
        SRAM_out_buffer[14]) );
  QDFFS window_reg_2__4__6_ ( .D(n3097), .CK(clk), .Q(window_2__4__6_) );
  QDFFS pool_temp_reg_1__6_ ( .D(n3078), .CK(clk), .Q(pool_temp[22]) );
  QDFFS pool_temp_reg_3__6_ ( .D(n3062), .CK(clk), .Q(pool_temp[6]) );
  QDFFS SRAM_out_buffer_reg_1__1__6_ ( .D(n3022), .CK(clk), .Q(
        SRAM_out_buffer[54]) );
  QDFFS SRAM_out_buffer_reg_0__1__6_ ( .D(n3021), .CK(clk), .Q(
        SRAM_out_buffer[86]) );
  QDFFS window_reg_1__3__6_ ( .D(n3020), .CK(clk), .Q(window_1__3__6_) );
  QDFFS window_reg_0__3__6_ ( .D(n3019), .CK(clk), .Q(window_0__3__6_) );
  QDFFS window_reg_1__1__6_ ( .D(n2935), .CK(clk), .Q(median_in[38]) );
  QDFFS window_reg_1__0__6_ ( .D(n2934), .CK(clk), .Q(median_in[46]) );
  QDFFS window_reg_0__2__6_ ( .D(n2933), .CK(clk), .Q(median_in[54]) );
  QDFFS window_reg_0__1__6_ ( .D(n2932), .CK(clk), .Q(median_in[62]) );
  QDFFS window_reg_0__0__6_ ( .D(n2931), .CK(clk), .Q(median_in[70]) );
  QDFFS SRAM_out_buffer_reg_2__1__6_ ( .D(n3018), .CK(clk), .Q(
        SRAM_out_buffer[22]) );
  QDFFS window_reg_2__3__6_ ( .D(n3017), .CK(clk), .Q(window_2__3__6_) );
  QDFFS window_reg_2__1__6_ ( .D(n2928), .CK(clk), .Q(median_in[14]) );
  QDFFS window_reg_2__0__6_ ( .D(n2927), .CK(clk), .Q(median_in[22]) );
  QDFFS filter_result_reg_reg_0__3__6_ ( .D(n3171), .CK(clk), .Q(
        filter_result_reg[70]) );
  QDFFS SRAM_64X32_data_in_reg_reg_6_ ( .D(n3061), .CK(clk), .Q(
        SRAM_64X32_in_decode[6]) );
  QDFFS filter_result_reg_reg_0__2__6_ ( .D(n3170), .CK(clk), .Q(
        filter_result_reg[78]) );
  QDFFS filter_result_reg_reg_0__1__6_ ( .D(n3169), .CK(clk), .Q(
        filter_result_reg[86]) );
  QDFFS SRAM_64X32_data_in_reg_reg_22_ ( .D(n3077), .CK(clk), .Q(
        SRAM_64X32_in_decode[22]) );
  QDFFS filter_result_reg_reg_0__0__6_ ( .D(n3168), .CK(clk), .Q(
        filter_result_reg[94]) );
  QDFFS pool_temp_reg_0__6_ ( .D(n2905), .CK(clk), .Q(pool_temp[30]) );
  QDFFS SRAM_64X32_data_in_reg_reg_30_ ( .D(n2904), .CK(clk), .Q(
        SRAM_64X32_in_decode[30]) );
  QDFFS pool_temp_reg_2__6_ ( .D(n2889), .CK(clk), .Q(pool_temp[14]) );
  QDFFS SRAM_64X32_data_in_reg_reg_14_ ( .D(n2888), .CK(clk), .Q(
        SRAM_64X32_in_decode[14]) );
  QDFFS SRAM_out_buffer_reg_1__2__5_ ( .D(n3108), .CK(clk), .Q(
        SRAM_out_buffer[45]) );
  QDFFS SRAM_out_buffer_reg_0__2__5_ ( .D(n3107), .CK(clk), .Q(
        SRAM_out_buffer[77]) );
  QDFFS window_reg_1__4__5_ ( .D(n3106), .CK(clk), .Q(window_1__4__5_) );
  QDFFS window_reg_0__4__5_ ( .D(n3105), .CK(clk), .Q(window_0__4__5_) );
  QDFFS SRAM_out_buffer_reg_2__2__5_ ( .D(n3104), .CK(clk), .Q(
        SRAM_out_buffer[13]) );
  QDFFS window_reg_2__4__5_ ( .D(n3103), .CK(clk), .Q(window_2__4__5_) );
  QDFFS pool_temp_reg_1__5_ ( .D(n3080), .CK(clk), .Q(pool_temp[21]) );
  QDFFS pool_temp_reg_3__5_ ( .D(n3064), .CK(clk), .Q(pool_temp[5]) );
  QDFFS SRAM_out_buffer_reg_1__1__5_ ( .D(n3028), .CK(clk), .Q(
        SRAM_out_buffer[53]) );
  QDFFS SRAM_out_buffer_reg_0__1__5_ ( .D(n3027), .CK(clk), .Q(
        SRAM_out_buffer[85]) );
  QDFFS window_reg_1__3__5_ ( .D(n3026), .CK(clk), .Q(window_1__3__5_) );
  QDFFS window_reg_0__3__5_ ( .D(n3025), .CK(clk), .Q(window_0__3__5_) );
  QDFFS window_reg_1__2__5_ ( .D(n2948), .CK(clk), .Q(median_in[29]) );
  QDFFS window_reg_1__1__5_ ( .D(n2947), .CK(clk), .Q(median_in[37]) );
  QDFFS window_reg_1__0__5_ ( .D(n2946), .CK(clk), .Q(median_in[45]) );
  QDFFS window_reg_0__1__5_ ( .D(n2944), .CK(clk), .Q(median_in[61]) );
  QDFFS window_reg_0__0__5_ ( .D(n2943), .CK(clk), .Q(median_in[69]) );
  QDFFS SRAM_out_buffer_reg_2__1__5_ ( .D(n3024), .CK(clk), .Q(
        SRAM_out_buffer[21]) );
  QDFFS window_reg_2__3__5_ ( .D(n3023), .CK(clk), .Q(window_2__3__5_) );
  QDFFS window_reg_2__2__5_ ( .D(n2941), .CK(clk), .Q(median_in[5]) );
  QDFFS window_reg_2__1__5_ ( .D(n2940), .CK(clk), .Q(median_in[13]) );
  QDFFS window_reg_2__0__5_ ( .D(n2939), .CK(clk), .Q(median_in[21]) );
  QDFFS filter_result_reg_reg_0__3__5_ ( .D(n3175), .CK(clk), .Q(
        filter_result_reg[69]) );
  QDFFS SRAM_64X32_data_in_reg_reg_5_ ( .D(n3063), .CK(clk), .Q(
        SRAM_64X32_in_decode[5]) );
  QDFFS filter_result_reg_reg_0__2__5_ ( .D(n3174), .CK(clk), .Q(
        filter_result_reg[77]) );
  QDFFS filter_result_reg_reg_0__1__5_ ( .D(n3173), .CK(clk), .Q(
        filter_result_reg[85]) );
  QDFFS SRAM_64X32_data_in_reg_reg_21_ ( .D(n3079), .CK(clk), .Q(
        SRAM_64X32_in_decode[21]) );
  QDFFS filter_result_reg_reg_0__0__5_ ( .D(n3172), .CK(clk), .Q(
        filter_result_reg[93]) );
  QDFFS pool_temp_reg_0__5_ ( .D(n2907), .CK(clk), .Q(pool_temp[29]) );
  QDFFS SRAM_64X32_data_in_reg_reg_29_ ( .D(n2906), .CK(clk), .Q(
        SRAM_64X32_in_decode[29]) );
  QDFFS pool_temp_reg_2__5_ ( .D(n2891), .CK(clk), .Q(pool_temp[13]) );
  QDFFS SRAM_64X32_data_in_reg_reg_13_ ( .D(n2890), .CK(clk), .Q(
        SRAM_64X32_in_decode[13]) );
  QDFFS SRAM_out_buffer_reg_1__2__4_ ( .D(n3114), .CK(clk), .Q(
        SRAM_out_buffer[44]) );
  QDFFS SRAM_out_buffer_reg_0__2__4_ ( .D(n3113), .CK(clk), .Q(
        SRAM_out_buffer[76]) );
  QDFFS window_reg_1__4__4_ ( .D(n3112), .CK(clk), .Q(window_1__4__4_) );
  QDFFS window_reg_0__4__4_ ( .D(n3111), .CK(clk), .Q(window_0__4__4_) );
  QDFFS SRAM_out_buffer_reg_2__2__4_ ( .D(n3110), .CK(clk), .Q(
        SRAM_out_buffer[12]) );
  QDFFS window_reg_2__4__4_ ( .D(n3109), .CK(clk), .Q(window_2__4__4_) );
  QDFFS pool_temp_reg_1__4_ ( .D(n3082), .CK(clk), .Q(pool_temp[20]) );
  QDFFS pool_temp_reg_3__4_ ( .D(n3066), .CK(clk), .Q(pool_temp[4]) );
  QDFFS SRAM_out_buffer_reg_1__1__4_ ( .D(n3034), .CK(clk), .Q(
        SRAM_out_buffer[52]) );
  QDFFS SRAM_out_buffer_reg_0__1__4_ ( .D(n3033), .CK(clk), .Q(
        SRAM_out_buffer[84]) );
  QDFFS window_reg_1__3__4_ ( .D(n3032), .CK(clk), .Q(window_1__3__4_) );
  QDFFS window_reg_0__3__4_ ( .D(n3031), .CK(clk), .Q(window_0__3__4_) );
  QDFFS window_reg_1__1__4_ ( .D(n2959), .CK(clk), .Q(median_in[36]) );
  QDFFS window_reg_1__0__4_ ( .D(n2958), .CK(clk), .Q(median_in[44]) );
  QDFFS window_reg_0__2__4_ ( .D(n2957), .CK(clk), .Q(median_in[52]) );
  QDFFS window_reg_0__1__4_ ( .D(n2956), .CK(clk), .Q(median_in[60]) );
  QDFFS window_reg_0__0__4_ ( .D(n2955), .CK(clk), .Q(median_in[68]) );
  QDFFS SRAM_out_buffer_reg_2__1__4_ ( .D(n3030), .CK(clk), .Q(
        SRAM_out_buffer[20]) );
  QDFFS window_reg_2__3__4_ ( .D(n3029), .CK(clk), .Q(window_2__3__4_) );
  QDFFS window_reg_2__1__4_ ( .D(n2952), .CK(clk), .Q(median_in[12]) );
  QDFFS window_reg_2__0__4_ ( .D(n2951), .CK(clk), .Q(median_in[20]) );
  QDFFS filter_result_reg_reg_0__3__4_ ( .D(n3179), .CK(clk), .Q(
        filter_result_reg[68]) );
  QDFFS SRAM_64X32_data_in_reg_reg_4_ ( .D(n3065), .CK(clk), .Q(
        SRAM_64X32_in_decode[4]) );
  QDFFS filter_result_reg_reg_0__2__4_ ( .D(n3178), .CK(clk), .Q(
        filter_result_reg[76]) );
  QDFFS filter_result_reg_reg_0__1__4_ ( .D(n3177), .CK(clk), .Q(
        filter_result_reg[84]) );
  QDFFS SRAM_64X32_data_in_reg_reg_20_ ( .D(n3081), .CK(clk), .Q(
        SRAM_64X32_in_decode[20]) );
  QDFFS filter_result_reg_reg_0__0__4_ ( .D(n3176), .CK(clk), .Q(
        filter_result_reg[92]) );
  QDFFS pool_temp_reg_0__4_ ( .D(n2909), .CK(clk), .Q(pool_temp[28]) );
  QDFFS SRAM_64X32_data_in_reg_reg_28_ ( .D(n2908), .CK(clk), .Q(
        SRAM_64X32_in_decode[28]) );
  QDFFS pool_temp_reg_2__4_ ( .D(n2893), .CK(clk), .Q(pool_temp[12]) );
  QDFFS SRAM_64X32_data_in_reg_reg_12_ ( .D(n2892), .CK(clk), .Q(
        SRAM_64X32_in_decode[12]) );
  QDFFS SRAM_out_buffer_reg_1__2__3_ ( .D(n3120), .CK(clk), .Q(
        SRAM_out_buffer[43]) );
  QDFFS SRAM_out_buffer_reg_0__2__3_ ( .D(n3119), .CK(clk), .Q(
        SRAM_out_buffer[75]) );
  QDFFS window_reg_1__4__3_ ( .D(n3118), .CK(clk), .Q(window_1__4__3_) );
  QDFFS window_reg_0__4__3_ ( .D(n3117), .CK(clk), .Q(window_0__4__3_) );
  QDFFS SRAM_out_buffer_reg_2__2__3_ ( .D(n3116), .CK(clk), .Q(
        SRAM_out_buffer[11]) );
  QDFFS window_reg_2__4__3_ ( .D(n3115), .CK(clk), .Q(window_2__4__3_) );
  QDFFS pool_temp_reg_1__3_ ( .D(n3084), .CK(clk), .Q(pool_temp[19]) );
  QDFFS pool_temp_reg_3__3_ ( .D(n3068), .CK(clk), .Q(pool_temp[3]) );
  QDFFS SRAM_out_buffer_reg_1__1__3_ ( .D(n3040), .CK(clk), .Q(
        SRAM_out_buffer[51]) );
  QDFFS SRAM_out_buffer_reg_0__1__3_ ( .D(n3039), .CK(clk), .Q(
        SRAM_out_buffer[83]) );
  QDFFS window_reg_1__3__3_ ( .D(n3038), .CK(clk), .Q(window_1__3__3_) );
  QDFFS window_reg_0__3__3_ ( .D(n3037), .CK(clk), .Q(window_0__3__3_) );
  QDFFS window_reg_1__1__3_ ( .D(n2971), .CK(clk), .Q(median_in[35]) );
  QDFFS window_reg_1__0__3_ ( .D(n2970), .CK(clk), .Q(median_in[43]) );
  QDFFS window_reg_0__2__3_ ( .D(n2969), .CK(clk), .Q(median_in[51]) );
  QDFFS window_reg_0__1__3_ ( .D(n2968), .CK(clk), .Q(median_in[59]) );
  QDFFS window_reg_0__0__3_ ( .D(n2967), .CK(clk), .Q(median_in[67]) );
  QDFFS SRAM_out_buffer_reg_2__1__3_ ( .D(n3036), .CK(clk), .Q(
        SRAM_out_buffer[19]) );
  QDFFS window_reg_2__3__3_ ( .D(n3035), .CK(clk), .Q(window_2__3__3_) );
  QDFFS window_reg_2__1__3_ ( .D(n2964), .CK(clk), .Q(median_in[11]) );
  QDFFS window_reg_2__0__3_ ( .D(n2963), .CK(clk), .Q(median_in[19]) );
  QDFFS filter_result_reg_reg_0__3__3_ ( .D(n3183), .CK(clk), .Q(
        filter_result_reg[67]) );
  QDFFS SRAM_64X32_data_in_reg_reg_3_ ( .D(n3067), .CK(clk), .Q(
        SRAM_64X32_in_decode[3]) );
  QDFFS filter_result_reg_reg_0__2__3_ ( .D(n3182), .CK(clk), .Q(
        filter_result_reg[75]) );
  QDFFS filter_result_reg_reg_0__1__3_ ( .D(n3181), .CK(clk), .Q(
        filter_result_reg[83]) );
  QDFFS SRAM_64X32_data_in_reg_reg_19_ ( .D(n3083), .CK(clk), .Q(
        SRAM_64X32_in_decode[19]) );
  QDFFS filter_result_reg_reg_0__0__3_ ( .D(n3180), .CK(clk), .Q(
        filter_result_reg[91]) );
  QDFFS pool_temp_reg_0__3_ ( .D(n2911), .CK(clk), .Q(pool_temp[27]) );
  QDFFS SRAM_64X32_data_in_reg_reg_27_ ( .D(n2910), .CK(clk), .Q(
        SRAM_64X32_in_decode[27]) );
  QDFFS pool_temp_reg_2__3_ ( .D(n2895), .CK(clk), .Q(pool_temp[11]) );
  QDFFS SRAM_64X32_data_in_reg_reg_11_ ( .D(n2894), .CK(clk), .Q(
        SRAM_64X32_in_decode[11]) );
  QDFFS SRAM_out_buffer_reg_1__2__2_ ( .D(n3126), .CK(clk), .Q(
        SRAM_out_buffer[42]) );
  QDFFS SRAM_out_buffer_reg_0__2__2_ ( .D(n3125), .CK(clk), .Q(
        SRAM_out_buffer[74]) );
  QDFFS window_reg_1__4__2_ ( .D(n3124), .CK(clk), .Q(window_1__4__2_) );
  QDFFS window_reg_0__4__2_ ( .D(n3123), .CK(clk), .Q(window_0__4__2_) );
  QDFFS SRAM_out_buffer_reg_2__2__2_ ( .D(n3122), .CK(clk), .Q(
        SRAM_out_buffer[10]) );
  QDFFS window_reg_2__4__2_ ( .D(n3121), .CK(clk), .Q(window_2__4__2_) );
  QDFFS pool_temp_reg_1__2_ ( .D(n3086), .CK(clk), .Q(pool_temp[18]) );
  QDFFS pool_temp_reg_3__2_ ( .D(n3070), .CK(clk), .Q(pool_temp[2]) );
  QDFFS SRAM_out_buffer_reg_1__1__2_ ( .D(n3046), .CK(clk), .Q(
        SRAM_out_buffer[50]) );
  QDFFS SRAM_out_buffer_reg_0__1__2_ ( .D(n3045), .CK(clk), .Q(
        SRAM_out_buffer[82]) );
  QDFFS window_reg_1__3__2_ ( .D(n3044), .CK(clk), .Q(window_1__3__2_) );
  QDFFS window_reg_0__3__2_ ( .D(n3043), .CK(clk), .Q(window_0__3__2_) );
  QDFFS window_reg_1__1__2_ ( .D(n2983), .CK(clk), .Q(median_in[34]) );
  QDFFS window_reg_0__2__2_ ( .D(n2981), .CK(clk), .Q(median_in[50]) );
  QDFFS window_reg_0__1__2_ ( .D(n2980), .CK(clk), .Q(median_in[58]) );
  QDFFS window_reg_0__0__2_ ( .D(n2979), .CK(clk), .Q(median_in[66]) );
  QDFFS SRAM_out_buffer_reg_2__1__2_ ( .D(n3042), .CK(clk), .Q(
        SRAM_out_buffer[18]) );
  QDFFS window_reg_2__3__2_ ( .D(n3041), .CK(clk), .Q(window_2__3__2_) );
  QDFFS window_reg_2__1__2_ ( .D(n2976), .CK(clk), .Q(median_in[10]) );
  QDFFS window_reg_2__0__2_ ( .D(n2975), .CK(clk), .Q(median_in[18]) );
  QDFFS filter_result_reg_reg_0__3__2_ ( .D(n3187), .CK(clk), .Q(
        filter_result_reg[66]) );
  QDFFS SRAM_64X32_data_in_reg_reg_2_ ( .D(n3069), .CK(clk), .Q(
        SRAM_64X32_in_decode[2]) );
  QDFFS filter_result_reg_reg_0__2__2_ ( .D(n3186), .CK(clk), .Q(
        filter_result_reg[74]) );
  QDFFS filter_result_reg_reg_0__1__2_ ( .D(n3185), .CK(clk), .Q(
        filter_result_reg[82]) );
  QDFFS SRAM_64X32_data_in_reg_reg_18_ ( .D(n3085), .CK(clk), .Q(
        SRAM_64X32_in_decode[18]) );
  QDFFS filter_result_reg_reg_0__0__2_ ( .D(n3184), .CK(clk), .Q(
        filter_result_reg[90]) );
  QDFFS pool_temp_reg_0__2_ ( .D(n2913), .CK(clk), .Q(pool_temp[26]) );
  QDFFS SRAM_64X32_data_in_reg_reg_26_ ( .D(n2912), .CK(clk), .Q(
        SRAM_64X32_in_decode[26]) );
  QDFFS pool_temp_reg_2__2_ ( .D(n2897), .CK(clk), .Q(pool_temp[10]) );
  QDFFS SRAM_64X32_data_in_reg_reg_10_ ( .D(n2896), .CK(clk), .Q(
        SRAM_64X32_in_decode[10]) );
  QDFFS SRAM_out_buffer_reg_1__3__1_ ( .D(n3159), .CK(clk), .Q(
        SRAM_out_buffer[33]) );
  QDFFS SRAM_out_buffer_reg_0__3__1_ ( .D(n3158), .CK(clk), .Q(
        SRAM_out_buffer[65]) );
  QDFFS window_reg_1__4__1_ ( .D(n3130), .CK(clk), .Q(window_1__4__1_) );
  QDFFS window_reg_1__3__1_ ( .D(n3050), .CK(clk), .Q(window_1__3__1_) );
  QDFFS window_reg_0__4__1_ ( .D(n3129), .CK(clk), .Q(window_0__4__1_) );
  QDFFS window_reg_0__3__1_ ( .D(n3049), .CK(clk), .Q(window_0__3__1_) );
  QDFFS SRAM_out_buffer_reg_2__3__1_ ( .D(n3157), .CK(clk), .Q(
        SRAM_out_buffer[1]) );
  QDFFS window_reg_2__4__1_ ( .D(n3127), .CK(clk), .Q(window_2__4__1_) );
  QDFFS window_reg_2__3__1_ ( .D(n3047), .CK(clk), .Q(window_2__3__1_) );
  QDFFS pool_temp_reg_1__1_ ( .D(n3088), .CK(clk), .Q(pool_temp[17]) );
  QDFFS pool_temp_reg_3__1_ ( .D(n3072), .CK(clk), .Q(pool_temp[1]) );
  QDFFS SRAM_out_buffer_reg_1__0__1_ ( .D(n2998), .CK(clk), .Q(
        SRAM_out_buffer[57]) );
  QDFFS SRAM_out_buffer_reg_0__0__1_ ( .D(n2997), .CK(clk), .Q(
        SRAM_out_buffer[89]) );
  QDFFS window_reg_1__1__1_ ( .D(n2995), .CK(clk), .Q(median_in[33]) );
  QDFFS window_reg_1__0__1_ ( .D(n2994), .CK(clk), .Q(median_in[41]) );
  QDFFS window_reg_0__2__1_ ( .D(n2993), .CK(clk), .Q(median_in[49]) );
  QDFFS window_reg_0__1__1_ ( .D(n2992), .CK(clk), .Q(median_in[57]) );
  QDFFS window_reg_0__0__1_ ( .D(n2991), .CK(clk), .Q(median_in[65]) );
  QDFFS SRAM_out_buffer_reg_2__0__1_ ( .D(n2990), .CK(clk), .Q(
        SRAM_out_buffer[25]) );
  QDFFS window_reg_2__1__1_ ( .D(n2988), .CK(clk), .Q(median_in[9]) );
  QDFFS window_reg_2__0__1_ ( .D(n2987), .CK(clk), .Q(median_in[17]) );
  QDFFS filter_result_reg_reg_0__3__1_ ( .D(n3191), .CK(clk), .Q(
        filter_result_reg[65]) );
  QDFFS SRAM_64X32_data_in_reg_reg_1_ ( .D(n3071), .CK(clk), .Q(
        SRAM_64X32_in_decode[1]) );
  QDFFS filter_result_reg_reg_0__2__1_ ( .D(n3190), .CK(clk), .Q(
        filter_result_reg[73]) );
  QDFFS filter_result_reg_reg_0__1__1_ ( .D(n3189), .CK(clk), .Q(
        filter_result_reg[81]) );
  QDFFS SRAM_64X32_data_in_reg_reg_17_ ( .D(n3087), .CK(clk), .Q(
        SRAM_64X32_in_decode[17]) );
  QDFFS filter_result_reg_reg_0__0__1_ ( .D(n3188), .CK(clk), .Q(
        filter_result_reg[89]) );
  QDFFS pool_temp_reg_0__1_ ( .D(n2915), .CK(clk), .Q(pool_temp[25]) );
  QDFFS SRAM_64X32_data_in_reg_reg_25_ ( .D(n2914), .CK(clk), .Q(
        SRAM_64X32_in_decode[25]) );
  QDFFS pool_temp_reg_2__1_ ( .D(n2899), .CK(clk), .Q(pool_temp[9]) );
  QDFFS SRAM_64X32_data_in_reg_reg_9_ ( .D(n2898), .CK(clk), .Q(
        SRAM_64X32_in_decode[9]) );
  QDFFS SRAM_out_buffer_reg_1__3__0_ ( .D(n3162), .CK(clk), .Q(
        SRAM_out_buffer[32]) );
  QDFFS SRAM_out_buffer_reg_0__3__0_ ( .D(n3161), .CK(clk), .Q(
        SRAM_out_buffer[64]) );
  QDFFS window_reg_1__4__0_ ( .D(n3136), .CK(clk), .Q(window_1__4__0_) );
  QDFFS window_reg_1__3__0_ ( .D(n3056), .CK(clk), .Q(window_1__3__0_) );
  QDFFS window_reg_0__4__0_ ( .D(n3135), .CK(clk), .Q(window_0__4__0_) );
  QDFFS window_reg_0__3__0_ ( .D(n3055), .CK(clk), .Q(window_0__3__0_) );
  QDFFS SRAM_out_buffer_reg_2__3__0_ ( .D(n3160), .CK(clk), .Q(
        SRAM_out_buffer[0]) );
  QDFFS window_reg_2__4__0_ ( .D(n3133), .CK(clk), .Q(window_2__4__0_) );
  QDFFS window_reg_2__3__0_ ( .D(n3053), .CK(clk), .Q(window_2__3__0_) );
  QDFFS pool_temp_reg_1__0_ ( .D(n3090), .CK(clk), .Q(pool_temp[16]) );
  QDFFS pool_temp_reg_3__0_ ( .D(n3074), .CK(clk), .Q(pool_temp[0]) );
  QDFFS SRAM_out_buffer_reg_1__0__0_ ( .D(n3010), .CK(clk), .Q(
        SRAM_out_buffer[56]) );
  QDFFS SRAM_out_buffer_reg_0__0__0_ ( .D(n3009), .CK(clk), .Q(
        SRAM_out_buffer[88]) );
  QDFFS window_reg_1__2__0_ ( .D(n3008), .CK(clk), .Q(median_in[24]) );
  QDFFS window_reg_1__1__0_ ( .D(n6305), .CK(clk), .Q(median_in[32]) );
  QDFFS window_reg_1__0__0_ ( .D(n3006), .CK(clk), .Q(median_in[40]) );
  QDFFS window_reg_0__1__0_ ( .D(n3004), .CK(clk), .Q(median_in[56]) );
  QDFFS window_reg_0__0__0_ ( .D(n3003), .CK(clk), .Q(median_in[64]) );
  QDFFS SRAM_out_buffer_reg_2__0__0_ ( .D(n3002), .CK(clk), .Q(
        SRAM_out_buffer[24]) );
  QDFFS window_reg_2__2__0_ ( .D(n3001), .CK(clk), .Q(median_in[0]) );
  QDFFS window_reg_2__1__0_ ( .D(n3000), .CK(clk), .Q(median_in[8]) );
  QDFFS window_reg_2__0__0_ ( .D(n2999), .CK(clk), .Q(median_in[16]) );
  QDFFS filter_result_reg_reg_0__3__0_ ( .D(n3195), .CK(clk), .Q(
        filter_result_reg[64]) );
  QDFFS SRAM_64X32_data_in_reg_reg_0_ ( .D(n3073), .CK(clk), .Q(
        SRAM_64X32_in_decode[0]) );
  QDFFS filter_result_reg_reg_0__2__0_ ( .D(n3194), .CK(clk), .Q(
        filter_result_reg[72]) );
  QDFFS filter_result_reg_reg_0__1__0_ ( .D(n3193), .CK(clk), .Q(
        filter_result_reg[80]) );
  QDFFS SRAM_64X32_data_in_reg_reg_16_ ( .D(n3089), .CK(clk), .Q(
        SRAM_64X32_in_decode[16]) );
  QDFFS filter_result_reg_reg_0__0__0_ ( .D(n3192), .CK(clk), .Q(
        filter_result_reg[88]) );
  QDFFS pool_temp_reg_0__0_ ( .D(n2917), .CK(clk), .Q(pool_temp[24]) );
  QDFFS SRAM_64X32_data_in_reg_reg_24_ ( .D(n2916), .CK(clk), .Q(
        SRAM_64X32_in_decode[24]) );
  QDFFS pool_temp_reg_2__0_ ( .D(n2901), .CK(clk), .Q(pool_temp[8]) );
  QDFFS SRAM_64X32_data_in_reg_reg_8_ ( .D(n2900), .CK(clk), .Q(
        SRAM_64X32_in_decode[8]) );
  QDFFRBS template_count_reg_0_ ( .D(n3343), .CK(clk), .RB(n6307), .Q(
        template_count[0]) );
  QDFFRBS template_count_reg_1_ ( .D(n3344), .CK(clk), .RB(n6306), .Q(
        template_count[1]) );
  QDFFRBS template_count_reg_2_ ( .D(n3345), .CK(clk), .RB(n6307), .Q(
        template_count[2]) );
  QDFFRBS template_count_reg_3_ ( .D(n3346), .CK(clk), .RB(n6307), .Q(
        template_count[3]) );
  QDFFRBS set_count_reg_0_ ( .D(n3400), .CK(clk), .RB(n3487), .Q(set_count[0])
         );
  QDFFRBS set_count_reg_1_ ( .D(n3197), .CK(clk), .RB(n6307), .Q(set_count[1])
         );
  QDFFRBS set_count_reg_2_ ( .D(n3399), .CK(clk), .RB(n6307), .Q(set_count[2])
         );
  QDFFRBS action_idx_reg_0_ ( .D(n3398), .CK(clk), .RB(n6307), .Q(
        action_idx[0]) );
  QDFFRBS action_idx_reg_1_ ( .D(n3397), .CK(clk), .RB(n6307), .Q(
        action_idx[1]) );
  QDFFRBS action_idx_reg_2_ ( .D(n3396), .CK(clk), .RB(n6307), .Q(
        action_idx[2]) );
  QDFFRBS action_idx_reg_3_ ( .D(n3395), .CK(clk), .RB(n6306), .Q(
        action_idx[3]) );
  QDFFRBS conv_dly3_reg_1_ ( .D(n3368), .CK(clk), .RB(n6307), .Q(conv_dly3[1])
         );
  QDFFRBS conv_dly3_reg_2_ ( .D(n3370), .CK(clk), .RB(n6306), .Q(conv_dly3[2])
         );
  QDFFRBS conv_dly3_reg_0_ ( .D(n3369), .CK(clk), .RB(n6307), .Q(conv_dly3[0])
         );
  QDFFRBS wait_conv_out_count_reg_3_ ( .D(n3363), .CK(clk), .RB(n6306), .Q(
        wait_conv_out_count[3]) );
  QDFFRBS wait_conv_out_count_reg_4_ ( .D(n3366), .CK(clk), .RB(n6307), .Q(
        wait_conv_out_count[4]) );
  QDFFRBS cal_count_reg_0_ ( .D(n3220), .CK(clk), .RB(n6306), .Q(cal_count[0])
         );
  QDFFRBS RGB_count_reg_0_ ( .D(N813), .CK(clk), .RB(n6307), .Q(RGB_count[0])
         );
  QDFFRBS RGB_count_reg_1_ ( .D(N814), .CK(clk), .RB(n6306), .Q(RGB_count[1])
         );
  QDFFRBS max_temp_reg_6_ ( .D(n3362), .CK(clk), .RB(n6307), .Q(max_temp[6])
         );
  QDFFRBS max_temp_reg_0_ ( .D(n3361), .CK(clk), .RB(n6307), .Q(max_temp[0])
         );
  QDFFRBS max_temp_reg_1_ ( .D(n3360), .CK(clk), .RB(n6307), .Q(max_temp[1])
         );
  QDFFRBS max_temp_reg_2_ ( .D(n3359), .CK(clk), .RB(n6307), .Q(max_temp[2])
         );
  QDFFRBS max_temp_reg_3_ ( .D(n3358), .CK(clk), .RB(n6307), .Q(max_temp[3])
         );
  QDFFRBS max_temp_reg_4_ ( .D(n3357), .CK(clk), .RB(n6307), .Q(max_temp[4])
         );
  QDFFRBS max_temp_reg_5_ ( .D(n3356), .CK(clk), .RB(n6307), .Q(max_temp[5])
         );
  QDFFRBS max_temp_reg_7_ ( .D(n3355), .CK(clk), .RB(n3487), .Q(max_temp[7])
         );
  QDFFRBS wgt_temp_reg_7_ ( .D(n3354), .CK(clk), .RB(n3487), .Q(wgt_temp[7])
         );
  QDFFRBS wgt_temp_reg_0_ ( .D(n3353), .CK(clk), .RB(n3487), .Q(wgt_temp[0])
         );
  QDFFRBS wgt_temp_reg_1_ ( .D(n3352), .CK(clk), .RB(n3487), .Q(wgt_temp[1])
         );
  QDFFRBS wgt_temp_reg_2_ ( .D(n3351), .CK(clk), .RB(n3487), .Q(wgt_temp[2])
         );
  QDFFRBS wgt_temp_reg_3_ ( .D(n3350), .CK(clk), .RB(n3487), .Q(wgt_temp[3])
         );
  QDFFRBS wgt_temp_reg_4_ ( .D(n3349), .CK(clk), .RB(n3487), .Q(wgt_temp[4])
         );
  QDFFRBS wgt_temp_reg_5_ ( .D(n3348), .CK(clk), .RB(n3487), .Q(wgt_temp[5])
         );
  QDFFRBS wgt_temp_reg_6_ ( .D(n3347), .CK(clk), .RB(n3487), .Q(wgt_temp[6])
         );
  QDFFRBS state_reg_1_ ( .D(n3404), .CK(clk), .RB(n3487), .Q(state[1]) );
  QDFFRBS SRAM_192_32_read_done_reg ( .D(n3229), .CK(clk), .RB(n3487), .Q(
        SRAM_192_32_read_done) );
  QDFFRBS cal_count_reg_8_ ( .D(n3235), .CK(clk), .RB(n6307), .Q(cal_count[8])
         );
  QDFFRBS cal_count_reg_5_ ( .D(n3225), .CK(clk), .RB(n6307), .Q(cal_count[5])
         );
  QDFFRBS cal_count_reg_4_ ( .D(n3224), .CK(clk), .RB(n6307), .Q(cal_count[4])
         );
  QDFFRBS SRAM_192_32_in_count_reg_0_ ( .D(n3269), .CK(clk), .RB(n6306), .Q(
        SRAM_192_32_in_count[0]) );
  QDFFRBS SRAM_192_32_in_count_reg_1_ ( .D(n3270), .CK(clk), .RB(n6306), .Q(
        SRAM_192_32_in_count[1]) );
  QDFFRBS start_write_flag_reg ( .D(n3268), .CK(clk), .RB(n6306), .Q(
        start_write_flag) );
  QDFFRBS SRAM_192X32_WE_reg ( .D(n6299), .CK(clk), .RB(n6306), .Q(
        SRAM_192X32_WE) );
  QDFFRBS cal_count_10_reg_0_ ( .D(n3217), .CK(clk), .RB(n6306), .Q(
        cal_count_10[0]) );
  QDFFRBS cal_count_10_reg_1_ ( .D(n3216), .CK(clk), .RB(n6306), .Q(
        cal_count_10[1]) );
  QDFFRBS cal_count_10_reg_2_ ( .D(n3218), .CK(clk), .RB(n6306), .Q(
        cal_count_10[2]) );
  QDFFRBS cal_count_10_reg_3_ ( .D(n3219), .CK(clk), .RB(n6306), .Q(
        cal_count_10[3]) );
  QDFFRBS cal_count_5_reg_0_ ( .D(n3215), .CK(clk), .RB(n6306), .Q(
        cal_count_5[0]) );
  QDFFRBS cal_count_5_reg_1_ ( .D(n3214), .CK(clk), .RB(n6306), .Q(
        cal_count_5[1]) );
  QDFFRBS cal_count_5_reg_2_ ( .D(n3213), .CK(clk), .RB(n6306), .Q(
        cal_count_5[2]) );
  QDFFRBS SRAM_64X32_WE_reg ( .D(n6300), .CK(clk), .RB(n6306), .Q(
        SRAM_64X32_WE) );
  QDFFRBS wb_addr_reg_7_ ( .D(n3205), .CK(clk), .RB(n6308), .Q(wb_addr[7]) );
  QDFFRBS wb_addr_reg_0_ ( .D(n3204), .CK(clk), .RB(n6308), .Q(wb_addr[0]) );
  QDFFRBS wb_addr_reg_1_ ( .D(n3203), .CK(clk), .RB(n3487), .Q(wb_addr[1]) );
  QDFFRBS wb_addr_reg_2_ ( .D(n3202), .CK(clk), .RB(n6308), .Q(wb_addr[2]) );
  QDFFRBS wb_addr_reg_3_ ( .D(n3201), .CK(clk), .RB(n6306), .Q(wb_addr[3]) );
  QDFFRBS wb_addr_reg_4_ ( .D(n3200), .CK(clk), .RB(n6308), .Q(wb_addr[4]) );
  QDFFRBS wb_addr_reg_5_ ( .D(n3199), .CK(clk), .RB(n6308), .Q(wb_addr[5]) );
  QDFFRBS wb_addr_reg_6_ ( .D(n3198), .CK(clk), .RB(n3487), .Q(wb_addr[6]) );
  QDFFRBS conv_temp_reg_1_ ( .D(n2882), .CK(clk), .RB(n6308), .Q(conv_temp[1])
         );
  QDFFRBS conv_temp_reg_2_ ( .D(n2881), .CK(clk), .RB(n6306), .Q(conv_temp[2])
         );
  QDFFRBS conv_temp_reg_3_ ( .D(n2880), .CK(clk), .RB(n6306), .Q(conv_temp[3])
         );
  QDFFRBS conv_temp_reg_4_ ( .D(n2879), .CK(clk), .RB(n6306), .Q(conv_temp[4])
         );
  QDFFRBS conv_temp_reg_5_ ( .D(n2878), .CK(clk), .RB(n6306), .Q(conv_temp[5])
         );
  QDFFRBS conv_temp_reg_6_ ( .D(n2877), .CK(clk), .RB(n6306), .Q(conv_temp[6])
         );
  QDFFRBS conv_temp_reg_7_ ( .D(n2876), .CK(clk), .RB(n6306), .Q(conv_temp[7])
         );
  QDFFRBS conv_temp_reg_8_ ( .D(n2875), .CK(clk), .RB(n6306), .Q(conv_temp[8])
         );
  QDFFRBS conv_temp_reg_9_ ( .D(n2874), .CK(clk), .RB(n6306), .Q(conv_temp[9])
         );
  QDFFRBS conv_temp_reg_10_ ( .D(n2873), .CK(clk), .RB(n6306), .Q(
        conv_temp[10]) );
  QDFFRBS conv_temp_reg_11_ ( .D(n2872), .CK(clk), .RB(n6306), .Q(
        conv_temp[11]) );
  QDFFRBS conv_temp_reg_12_ ( .D(n2871), .CK(clk), .RB(n6306), .Q(
        conv_temp[12]) );
  QDFFRBS conv_temp_reg_13_ ( .D(n2870), .CK(clk), .RB(n6306), .Q(
        conv_temp[13]) );
  QDFFRBS conv_temp_reg_14_ ( .D(n2869), .CK(clk), .RB(n6306), .Q(
        conv_temp[14]) );
  QDFFRBS conv_temp_reg_15_ ( .D(n2868), .CK(clk), .RB(n6306), .Q(
        conv_temp[15]) );
  QDFFRBS conv_temp_reg_16_ ( .D(n2867), .CK(clk), .RB(n6306), .Q(
        conv_temp[16]) );
  QDFFRBS conv_temp_reg_17_ ( .D(n2866), .CK(clk), .RB(n6306), .Q(
        conv_temp[17]) );
  QDFFRBS conv_temp_reg_18_ ( .D(n2865), .CK(clk), .RB(rst_n), .Q(
        conv_temp[18]) );
  QDFFRBS conv_temp_reg_19_ ( .D(n2862), .CK(clk), .RB(n6308), .Q(
        conv_temp[19]) );
  QDFFRBS find_median_inst_max3_reg_reg_7_ ( .D(find_median_inst_max3[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max3_reg[7]) );
  QDFFRBS find_median_inst_max_min_reg_reg_7_ ( .D(find_median_inst_max_min[7]), .CK(clk), .RB(n6308), .Q(find_median_inst_max_min_reg[7]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_7_ ( .D(
        find_median_inst_final_mid[7]), .CK(clk), .RB(n6308), .Q(
        median_result[7]) );
  QDFFRBS find_median_inst_mid2_reg_reg_7_ ( .D(find_median_inst_mid2[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid2_reg[7]) );
  QDFFRBS find_median_inst_min2_reg_reg_7_ ( .D(find_median_inst_min2[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min2_reg[7]) );
  QDFFRBS find_median_inst_max2_reg_reg_7_ ( .D(find_median_inst_max2[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max2_reg[7]) );
  QDFFRBS find_median_inst_mid1_reg_reg_7_ ( .D(find_median_inst_mid1[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid1_reg[7]) );
  QDFFRBS find_median_inst_min1_reg_reg_7_ ( .D(find_median_inst_min1[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min1_reg[7]) );
  QDFFRBS find_median_inst_max1_reg_reg_7_ ( .D(find_median_inst_max1[7]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max1_reg[7]) );
  QDFFRBS find_median_inst_mid3_reg_reg_7_ ( .D(find_median_inst_mid3[7]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid3_reg[7]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_7_ ( .D(find_median_inst_mid_mid[7]), .CK(clk), .RB(n3487), .Q(find_median_inst_mid_mid_reg[7]) );
  QDFFRBS find_median_inst_min3_reg_reg_7_ ( .D(find_median_inst_min3[7]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min3_reg[7]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_7_ ( .D(
        find_median_inst_min_max[7]), .CK(clk), .RB(n3487), .Q(
        find_median_inst_min_pool_temp[7]) );
  QDFFRBS find_median_inst_mid2_reg_reg_6_ ( .D(find_median_inst_mid2[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid2_reg[6]) );
  QDFFRBS find_median_inst_min2_reg_reg_6_ ( .D(find_median_inst_min2[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min2_reg[6]) );
  QDFFRBS find_median_inst_max2_reg_reg_6_ ( .D(find_median_inst_max2[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max2_reg[6]) );
  QDFFRBS find_median_inst_mid1_reg_reg_6_ ( .D(find_median_inst_mid1[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid1_reg[6]) );
  QDFFRBS find_median_inst_min1_reg_reg_6_ ( .D(find_median_inst_min1[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min1_reg[6]) );
  QDFFRBS find_median_inst_max1_reg_reg_6_ ( .D(find_median_inst_max1[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max1_reg[6]) );
  QDFFRBS find_median_inst_mid3_reg_reg_6_ ( .D(find_median_inst_mid3[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid3_reg[6]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_6_ ( .D(find_median_inst_mid_mid[6]), .CK(clk), .RB(n3487), .Q(find_median_inst_mid_mid_reg[6]) );
  QDFFRBS find_median_inst_min3_reg_reg_6_ ( .D(find_median_inst_min3[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min3_reg[6]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_6_ ( .D(
        find_median_inst_min_max[6]), .CK(clk), .RB(n3487), .Q(
        find_median_inst_min_pool_temp[6]) );
  QDFFRBS find_median_inst_max3_reg_reg_6_ ( .D(find_median_inst_max3[6]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max3_reg[6]) );
  QDFFRBS find_median_inst_max_min_reg_reg_6_ ( .D(find_median_inst_max_min[6]), .CK(clk), .RB(n3487), .Q(find_median_inst_max_min_reg[6]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_6_ ( .D(
        find_median_inst_final_mid[6]), .CK(clk), .RB(n3487), .Q(
        median_result[6]) );
  QDFFRBS find_median_inst_mid2_reg_reg_5_ ( .D(find_median_inst_mid2[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid2_reg[5]) );
  QDFFRBS find_median_inst_min2_reg_reg_5_ ( .D(find_median_inst_min2[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min2_reg[5]) );
  QDFFRBS find_median_inst_max2_reg_reg_5_ ( .D(find_median_inst_max2[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max2_reg[5]) );
  QDFFRBS find_median_inst_mid1_reg_reg_5_ ( .D(find_median_inst_mid1[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid1_reg[5]) );
  QDFFRBS find_median_inst_min1_reg_reg_5_ ( .D(find_median_inst_min1[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min1_reg[5]) );
  QDFFRBS find_median_inst_max1_reg_reg_5_ ( .D(find_median_inst_max1[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max1_reg[5]) );
  QDFFRBS find_median_inst_mid3_reg_reg_5_ ( .D(find_median_inst_mid3[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid3_reg[5]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_5_ ( .D(find_median_inst_mid_mid[5]), .CK(clk), .RB(n3487), .Q(find_median_inst_mid_mid_reg[5]) );
  QDFFRBS find_median_inst_min3_reg_reg_5_ ( .D(find_median_inst_min3[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min3_reg[5]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_5_ ( .D(
        find_median_inst_min_max[5]), .CK(clk), .RB(n3487), .Q(
        find_median_inst_min_pool_temp[5]) );
  QDFFRBS find_median_inst_max3_reg_reg_5_ ( .D(find_median_inst_max3[5]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max3_reg[5]) );
  QDFFRBS find_median_inst_max_min_reg_reg_5_ ( .D(find_median_inst_max_min[5]), .CK(clk), .RB(n3487), .Q(find_median_inst_max_min_reg[5]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_5_ ( .D(
        find_median_inst_final_mid[5]), .CK(clk), .RB(n3487), .Q(
        median_result[5]) );
  QDFFRBS find_median_inst_mid2_reg_reg_4_ ( .D(find_median_inst_mid2[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid2_reg[4]) );
  QDFFRBS find_median_inst_min2_reg_reg_4_ ( .D(find_median_inst_min2[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min2_reg[4]) );
  QDFFRBS find_median_inst_max2_reg_reg_4_ ( .D(find_median_inst_max2[4]), 
        .CK(clk), .RB(rst_n), .Q(find_median_inst_max2_reg[4]) );
  QDFFRBS find_median_inst_mid1_reg_reg_4_ ( .D(find_median_inst_mid1[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid1_reg[4]) );
  QDFFRBS find_median_inst_min1_reg_reg_4_ ( .D(find_median_inst_min1[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min1_reg[4]) );
  QDFFRBS find_median_inst_max1_reg_reg_4_ ( .D(find_median_inst_max1[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max1_reg[4]) );
  QDFFRBS find_median_inst_mid3_reg_reg_4_ ( .D(find_median_inst_mid3[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid3_reg[4]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_4_ ( .D(find_median_inst_mid_mid[4]), .CK(clk), .RB(n3487), .Q(find_median_inst_mid_mid_reg[4]) );
  QDFFRBS find_median_inst_min3_reg_reg_4_ ( .D(find_median_inst_min3[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min3_reg[4]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_4_ ( .D(
        find_median_inst_min_max[4]), .CK(clk), .RB(n3487), .Q(
        find_median_inst_min_pool_temp[4]) );
  QDFFRBS find_median_inst_max3_reg_reg_4_ ( .D(find_median_inst_max3[4]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max3_reg[4]) );
  QDFFRBS find_median_inst_max_min_reg_reg_4_ ( .D(find_median_inst_max_min[4]), .CK(clk), .RB(n3487), .Q(find_median_inst_max_min_reg[4]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_4_ ( .D(
        find_median_inst_final_mid[4]), .CK(clk), .RB(n3487), .Q(
        median_result[4]) );
  QDFFRBS find_median_inst_mid2_reg_reg_3_ ( .D(find_median_inst_mid2[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid2_reg[3]) );
  QDFFRBS find_median_inst_min2_reg_reg_3_ ( .D(find_median_inst_min2[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min2_reg[3]) );
  QDFFRBS find_median_inst_max2_reg_reg_3_ ( .D(find_median_inst_max2[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max2_reg[3]) );
  QDFFRBS find_median_inst_mid1_reg_reg_3_ ( .D(find_median_inst_mid1[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid1_reg[3]) );
  QDFFRBS find_median_inst_min1_reg_reg_3_ ( .D(find_median_inst_min1[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min1_reg[3]) );
  QDFFRBS find_median_inst_max1_reg_reg_3_ ( .D(find_median_inst_max1[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max1_reg[3]) );
  QDFFRBS find_median_inst_mid3_reg_reg_3_ ( .D(find_median_inst_mid3[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_mid3_reg[3]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_3_ ( .D(find_median_inst_mid_mid[3]), .CK(clk), .RB(n3487), .Q(find_median_inst_mid_mid_reg[3]) );
  QDFFRBS find_median_inst_min3_reg_reg_3_ ( .D(find_median_inst_min3[3]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_min3_reg[3]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_3_ ( .D(
        find_median_inst_min_max[3]), .CK(clk), .RB(n6308), .Q(
        find_median_inst_min_pool_temp[3]) );
  QDFFRBS find_median_inst_max3_reg_reg_3_ ( .D(find_median_inst_max3[3]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max3_reg[3]) );
  QDFFRBS find_median_inst_max_min_reg_reg_3_ ( .D(find_median_inst_max_min[3]), .CK(clk), .RB(n6308), .Q(find_median_inst_max_min_reg[3]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_3_ ( .D(
        find_median_inst_final_mid[3]), .CK(clk), .RB(n6308), .Q(
        median_result[3]) );
  QDFFRBS find_median_inst_mid2_reg_reg_2_ ( .D(find_median_inst_mid2[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid2_reg[2]) );
  QDFFRBS find_median_inst_min2_reg_reg_2_ ( .D(find_median_inst_min2[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min2_reg[2]) );
  QDFFRBS find_median_inst_max2_reg_reg_2_ ( .D(find_median_inst_max2[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max2_reg[2]) );
  QDFFRBS find_median_inst_mid1_reg_reg_2_ ( .D(find_median_inst_mid1[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid1_reg[2]) );
  QDFFRBS find_median_inst_min1_reg_reg_2_ ( .D(find_median_inst_min1[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min1_reg[2]) );
  QDFFRBS find_median_inst_max1_reg_reg_2_ ( .D(find_median_inst_max1[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max1_reg[2]) );
  QDFFRBS find_median_inst_mid3_reg_reg_2_ ( .D(find_median_inst_mid3[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid3_reg[2]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_2_ ( .D(find_median_inst_mid_mid[2]), .CK(clk), .RB(n6308), .Q(find_median_inst_mid_mid_reg[2]) );
  QDFFRBS find_median_inst_min3_reg_reg_2_ ( .D(find_median_inst_min3[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min3_reg[2]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_2_ ( .D(
        find_median_inst_min_max[2]), .CK(clk), .RB(n6308), .Q(
        find_median_inst_min_pool_temp[2]) );
  QDFFRBS find_median_inst_max3_reg_reg_2_ ( .D(find_median_inst_max3[2]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max3_reg[2]) );
  QDFFRBS find_median_inst_max_min_reg_reg_2_ ( .D(find_median_inst_max_min[2]), .CK(clk), .RB(n6308), .Q(find_median_inst_max_min_reg[2]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_2_ ( .D(
        find_median_inst_final_mid[2]), .CK(clk), .RB(n6308), .Q(
        median_result[2]) );
  QDFFRBS find_median_inst_mid2_reg_reg_1_ ( .D(find_median_inst_mid2[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid2_reg[1]) );
  QDFFRBS find_median_inst_max2_reg_reg_1_ ( .D(find_median_inst_max2[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max2_reg[1]) );
  QDFFRBS find_median_inst_mid1_reg_reg_1_ ( .D(find_median_inst_mid1[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid1_reg[1]) );
  QDFFRBS find_median_inst_mid3_reg_reg_1_ ( .D(find_median_inst_mid3[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid3_reg[1]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_1_ ( .D(find_median_inst_mid_mid[1]), .CK(clk), .RB(n6308), .Q(find_median_inst_mid_mid_reg[1]) );
  QDFFRBS find_median_inst_min3_reg_reg_1_ ( .D(find_median_inst_min3[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min3_reg[1]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_1_ ( .D(
        find_median_inst_min_max[1]), .CK(clk), .RB(n6308), .Q(
        find_median_inst_min_pool_temp[1]) );
  QDFFRBS find_median_inst_max3_reg_reg_1_ ( .D(find_median_inst_max3[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max3_reg[1]) );
  QDFFRBS find_median_inst_max_min_reg_reg_1_ ( .D(find_median_inst_max_min[1]), .CK(clk), .RB(n6308), .Q(find_median_inst_max_min_reg[1]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_1_ ( .D(
        find_median_inst_final_mid[1]), .CK(clk), .RB(n6308), .Q(
        median_result[1]) );
  QDFFRBS find_median_inst_mid2_reg_reg_0_ ( .D(find_median_inst_mid2[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid2_reg[0]) );
  QDFFRBS find_median_inst_min2_reg_reg_0_ ( .D(find_median_inst_min2[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min2_reg[0]) );
  QDFFRBS find_median_inst_max2_reg_reg_0_ ( .D(find_median_inst_max2[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max2_reg[0]) );
  QDFFRBS find_median_inst_mid1_reg_reg_0_ ( .D(find_median_inst_mid1[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid1_reg[0]) );
  QDFFRBS find_median_inst_max1_reg_reg_0_ ( .D(find_median_inst_max1[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max1_reg[0]) );
  QDFFRBS find_median_inst_mid3_reg_reg_0_ ( .D(find_median_inst_mid3[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_mid3_reg[0]) );
  QDFFRBS find_median_inst_mid_mid_reg_reg_0_ ( .D(find_median_inst_mid_mid[0]), .CK(clk), .RB(n6308), .Q(find_median_inst_mid_mid_reg[0]) );
  QDFFRBS find_median_inst_min3_reg_reg_0_ ( .D(find_median_inst_min3[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min3_reg[0]) );
  QDFFRBS find_median_inst_min_pool_temp_reg_0_ ( .D(
        find_median_inst_min_max[0]), .CK(clk), .RB(n6308), .Q(
        find_median_inst_min_pool_temp[0]) );
  QDFFRBS find_median_inst_max3_reg_reg_0_ ( .D(find_median_inst_max3[0]), 
        .CK(clk), .RB(n3487), .Q(find_median_inst_max3_reg[0]) );
  QDFFRBS find_median_inst_max_min_reg_reg_0_ ( .D(find_median_inst_max_min[0]), .CK(clk), .RB(rst_n), .Q(find_median_inst_max_min_reg[0]) );
  QDFFRBS find_median_inst_final_mid_reg_reg_0_ ( .D(
        find_median_inst_final_mid[0]), .CK(clk), .RB(n6308), .Q(
        median_result[0]) );
  QDFFS image_size_reg_reg_0_ ( .D(n2861), .CK(clk), .Q(image_size_reg[0]) );
  QDFFS image_size_reg_reg_1_ ( .D(n2860), .CK(clk), .Q(image_size_reg[1]) );
  QDFFS conv_out_reg_reg_0_ ( .D(n2859), .CK(clk), .Q(conv_out_reg[0]) );
  QDFFS conv_out_reg_reg_19_ ( .D(n2858), .CK(clk), .Q(conv_out_reg[19]) );
  QDFFS conv_out_reg_reg_18_ ( .D(n2857), .CK(clk), .Q(conv_out_reg[18]) );
  QDFFS conv_out_reg_reg_17_ ( .D(n2856), .CK(clk), .Q(conv_out_reg[17]) );
  QDFFS conv_out_reg_reg_16_ ( .D(n2855), .CK(clk), .Q(conv_out_reg[16]) );
  QDFFS conv_out_reg_reg_15_ ( .D(n2854), .CK(clk), .Q(conv_out_reg[15]) );
  QDFFS conv_out_reg_reg_14_ ( .D(n2853), .CK(clk), .Q(conv_out_reg[14]) );
  QDFFS conv_out_reg_reg_13_ ( .D(n2852), .CK(clk), .Q(conv_out_reg[13]) );
  QDFFS conv_out_reg_reg_12_ ( .D(n2851), .CK(clk), .Q(conv_out_reg[12]) );
  QDFFS conv_out_reg_reg_11_ ( .D(n2850), .CK(clk), .Q(conv_out_reg[11]) );
  QDFFS conv_out_reg_reg_10_ ( .D(n2849), .CK(clk), .Q(conv_out_reg[10]) );
  QDFFS conv_out_reg_reg_9_ ( .D(n2848), .CK(clk), .Q(conv_out_reg[9]) );
  QDFFS conv_out_reg_reg_8_ ( .D(n2847), .CK(clk), .Q(conv_out_reg[8]) );
  QDFFS conv_out_reg_reg_7_ ( .D(n2846), .CK(clk), .Q(conv_out_reg[7]) );
  QDFFS conv_out_reg_reg_6_ ( .D(n2845), .CK(clk), .Q(conv_out_reg[6]) );
  QDFFS conv_out_reg_reg_5_ ( .D(n2844), .CK(clk), .Q(conv_out_reg[5]) );
  QDFFS conv_out_reg_reg_4_ ( .D(n2843), .CK(clk), .Q(conv_out_reg[4]) );
  QDFFS conv_out_reg_reg_3_ ( .D(n2842), .CK(clk), .Q(conv_out_reg[3]) );
  QDFFS conv_out_reg_reg_2_ ( .D(n2841), .CK(clk), .Q(conv_out_reg[2]) );
  QDFFS conv_out_reg_reg_1_ ( .D(n2840), .CK(clk), .Q(conv_out_reg[1]) );
  QDFFS gray_wgt_reg_reg_0__7_ ( .D(n2839), .CK(clk), .Q(gray_wgt_reg[31]) );
  QDFFS gray_wgt_reg_reg_0__6_ ( .D(n2838), .CK(clk), .Q(gray_wgt_reg[30]) );
  QDFFS gray_wgt_reg_reg_0__5_ ( .D(n2837), .CK(clk), .Q(gray_wgt_reg[29]) );
  QDFFS gray_wgt_reg_reg_0__4_ ( .D(n2836), .CK(clk), .Q(gray_wgt_reg[28]) );
  QDFFS gray_wgt_reg_reg_0__3_ ( .D(n2835), .CK(clk), .Q(gray_wgt_reg[27]) );
  QDFFS gray_wgt_reg_reg_0__2_ ( .D(n2834), .CK(clk), .Q(gray_wgt_reg[26]) );
  QDFFS gray_wgt_reg_reg_0__1_ ( .D(n2833), .CK(clk), .Q(gray_wgt_reg[25]) );
  QDFFS gray_wgt_reg_reg_0__0_ ( .D(n2832), .CK(clk), .Q(gray_wgt_reg[24]) );
  QDFFS gray_wgt_reg_reg_1__7_ ( .D(n2831), .CK(clk), .Q(gray_wgt_reg[23]) );
  QDFFS gray_wgt_reg_reg_1__6_ ( .D(n2830), .CK(clk), .Q(gray_wgt_reg[22]) );
  QDFFS gray_wgt_reg_reg_1__5_ ( .D(n2829), .CK(clk), .Q(gray_wgt_reg[21]) );
  QDFFS gray_wgt_reg_reg_1__4_ ( .D(n2828), .CK(clk), .Q(gray_wgt_reg[20]) );
  QDFFS gray_wgt_reg_reg_1__3_ ( .D(n2827), .CK(clk), .Q(gray_wgt_reg[19]) );
  QDFFS gray_wgt_reg_reg_1__2_ ( .D(n2826), .CK(clk), .Q(gray_wgt_reg[18]) );
  QDFFS gray_wgt_reg_reg_1__1_ ( .D(n2825), .CK(clk), .Q(gray_wgt_reg[17]) );
  QDFFS gray_wgt_reg_reg_1__0_ ( .D(n2824), .CK(clk), .Q(gray_wgt_reg[16]) );
  QDFFS gray_wgt_reg_reg_2__7_ ( .D(n2823), .CK(clk), .Q(gray_wgt_reg[15]) );
  QDFFS gray_wgt_reg_reg_2__6_ ( .D(n2822), .CK(clk), .Q(gray_wgt_reg[14]) );
  QDFFS gray_wgt_reg_reg_2__5_ ( .D(n2821), .CK(clk), .Q(gray_wgt_reg[13]) );
  QDFFS gray_wgt_reg_reg_2__4_ ( .D(n2820), .CK(clk), .Q(gray_wgt_reg[12]) );
  QDFFS gray_wgt_reg_reg_2__3_ ( .D(n2819), .CK(clk), .Q(gray_wgt_reg[11]) );
  QDFFS gray_wgt_reg_reg_2__2_ ( .D(n2818), .CK(clk), .Q(gray_wgt_reg[10]) );
  QDFFS gray_wgt_reg_reg_2__1_ ( .D(n2817), .CK(clk), .Q(gray_wgt_reg[9]) );
  QDFFS gray_wgt_reg_reg_2__0_ ( .D(n2816), .CK(clk), .Q(gray_wgt_reg[8]) );
  QDFFS gray_wgt_reg_reg_3__0_ ( .D(n2815), .CK(clk), .Q(gray_wgt_reg[0]) );
  QDFFS gray_wgt_reg_reg_3__7_ ( .D(n2814), .CK(clk), .Q(gray_wgt_reg[7]) );
  QDFFS gray_wgt_reg_reg_3__6_ ( .D(n2813), .CK(clk), .Q(gray_wgt_reg[6]) );
  QDFFS gray_wgt_reg_reg_3__5_ ( .D(n2812), .CK(clk), .Q(gray_wgt_reg[5]) );
  QDFFS gray_wgt_reg_reg_3__4_ ( .D(n2811), .CK(clk), .Q(gray_wgt_reg[4]) );
  QDFFS gray_wgt_reg_reg_3__3_ ( .D(n2810), .CK(clk), .Q(gray_wgt_reg[3]) );
  QDFFS gray_wgt_reg_reg_3__2_ ( .D(n2809), .CK(clk), .Q(gray_wgt_reg[2]) );
  QDFFS gray_wgt_reg_reg_3__1_ ( .D(n2808), .CK(clk), .Q(gray_wgt_reg[1]) );
  QDFFS gray_max_temp_reg_0__6_ ( .D(n2807), .CK(clk), .Q(gray_max_temp[30])
         );
  QDFFS gray_max_temp_reg_1__6_ ( .D(n2806), .CK(clk), .Q(gray_max_temp[22])
         );
  QDFFS gray_max_temp_reg_2__6_ ( .D(n2805), .CK(clk), .Q(gray_max_temp[14])
         );
  QDFFS gray_max_temp_reg_3__6_ ( .D(n2804), .CK(clk), .Q(gray_max_temp[6]) );
  QDFFS gray_max_temp_reg_0__0_ ( .D(n2803), .CK(clk), .Q(gray_max_temp[24])
         );
  QDFFS gray_max_temp_reg_1__0_ ( .D(n2802), .CK(clk), .Q(gray_max_temp[16])
         );
  QDFFS gray_max_temp_reg_2__0_ ( .D(n2801), .CK(clk), .Q(gray_max_temp[8]) );
  QDFFS gray_max_temp_reg_3__0_ ( .D(n2800), .CK(clk), .Q(gray_max_temp[0]) );
  QDFFS gray_max_temp_reg_0__1_ ( .D(n2799), .CK(clk), .Q(gray_max_temp[25])
         );
  QDFFS gray_max_temp_reg_1__1_ ( .D(n2798), .CK(clk), .Q(gray_max_temp[17])
         );
  QDFFS gray_max_temp_reg_2__1_ ( .D(n2797), .CK(clk), .Q(gray_max_temp[9]) );
  QDFFS gray_max_temp_reg_3__1_ ( .D(n2796), .CK(clk), .Q(gray_max_temp[1]) );
  QDFFS gray_max_temp_reg_0__2_ ( .D(n2795), .CK(clk), .Q(gray_max_temp[26])
         );
  QDFFS gray_max_temp_reg_1__2_ ( .D(n2794), .CK(clk), .Q(gray_max_temp[18])
         );
  QDFFS gray_max_temp_reg_2__2_ ( .D(n2793), .CK(clk), .Q(gray_max_temp[10])
         );
  QDFFS gray_max_temp_reg_3__2_ ( .D(n2792), .CK(clk), .Q(gray_max_temp[2]) );
  QDFFS gray_max_temp_reg_0__3_ ( .D(n2791), .CK(clk), .Q(gray_max_temp[27])
         );
  QDFFS gray_max_temp_reg_1__3_ ( .D(n2790), .CK(clk), .Q(gray_max_temp[19])
         );
  QDFFS gray_max_temp_reg_2__3_ ( .D(n2789), .CK(clk), .Q(gray_max_temp[11])
         );
  QDFFS gray_max_temp_reg_3__3_ ( .D(n2788), .CK(clk), .Q(gray_max_temp[3]) );
  QDFFS gray_max_temp_reg_0__4_ ( .D(n2787), .CK(clk), .Q(gray_max_temp[28])
         );
  QDFFS gray_max_temp_reg_1__4_ ( .D(n2786), .CK(clk), .Q(gray_max_temp[20])
         );
  QDFFS gray_max_temp_reg_2__4_ ( .D(n2785), .CK(clk), .Q(gray_max_temp[12])
         );
  QDFFS gray_max_temp_reg_3__4_ ( .D(n2784), .CK(clk), .Q(gray_max_temp[4]) );
  QDFFS gray_max_temp_reg_0__5_ ( .D(n2783), .CK(clk), .Q(gray_max_temp[29])
         );
  QDFFS gray_max_temp_reg_1__5_ ( .D(n2782), .CK(clk), .Q(gray_max_temp[21])
         );
  QDFFS gray_max_temp_reg_2__5_ ( .D(n2781), .CK(clk), .Q(gray_max_temp[13])
         );
  QDFFS gray_max_temp_reg_3__5_ ( .D(n2780), .CK(clk), .Q(gray_max_temp[5]) );
  QDFFS gray_max_temp_reg_0__7_ ( .D(n2779), .CK(clk), .Q(gray_max_temp[31])
         );
  QDFFS gray_max_temp_reg_1__7_ ( .D(n2778), .CK(clk), .Q(gray_max_temp[23])
         );
  QDFFS gray_max_temp_reg_2__7_ ( .D(n2777), .CK(clk), .Q(gray_max_temp[15])
         );
  QDFFS gray_max_temp_reg_3__7_ ( .D(n2776), .CK(clk), .Q(gray_max_temp[7]) );
  QDFFS gray_avg_reg_reg_0__7_ ( .D(n2775), .CK(clk), .Q(gray_avg_reg[31]) );
  QDFFS gray_avg_reg_reg_0__6_ ( .D(n2774), .CK(clk), .Q(gray_avg_reg[30]) );
  QDFFS gray_avg_reg_reg_0__5_ ( .D(n2773), .CK(clk), .Q(gray_avg_reg[29]) );
  QDFFS gray_avg_reg_reg_0__4_ ( .D(n2772), .CK(clk), .Q(gray_avg_reg[28]) );
  QDFFS gray_avg_reg_reg_0__3_ ( .D(n2771), .CK(clk), .Q(gray_avg_reg[27]) );
  QDFFS gray_avg_reg_reg_0__2_ ( .D(n2770), .CK(clk), .Q(gray_avg_reg[26]) );
  QDFFS gray_avg_reg_reg_0__1_ ( .D(n2769), .CK(clk), .Q(gray_avg_reg[25]) );
  QDFFS gray_avg_reg_reg_0__0_ ( .D(n2768), .CK(clk), .Q(gray_avg_reg[24]) );
  QDFFS gray_avg_reg_reg_1__7_ ( .D(n2767), .CK(clk), .Q(gray_avg_reg[23]) );
  QDFFS gray_avg_reg_reg_1__6_ ( .D(n2766), .CK(clk), .Q(gray_avg_reg[22]) );
  QDFFS gray_avg_reg_reg_1__5_ ( .D(n2765), .CK(clk), .Q(gray_avg_reg[21]) );
  QDFFS gray_avg_reg_reg_1__4_ ( .D(n2764), .CK(clk), .Q(gray_avg_reg[20]) );
  QDFFS gray_avg_reg_reg_1__3_ ( .D(n2763), .CK(clk), .Q(gray_avg_reg[19]) );
  QDFFS gray_avg_reg_reg_1__2_ ( .D(n2762), .CK(clk), .Q(gray_avg_reg[18]) );
  QDFFS gray_avg_reg_reg_1__1_ ( .D(n2761), .CK(clk), .Q(gray_avg_reg[17]) );
  QDFFS gray_avg_reg_reg_1__0_ ( .D(n2760), .CK(clk), .Q(gray_avg_reg[16]) );
  QDFFS gray_avg_reg_reg_2__7_ ( .D(n2759), .CK(clk), .Q(gray_avg_reg[15]) );
  QDFFS gray_avg_reg_reg_2__6_ ( .D(n2758), .CK(clk), .Q(gray_avg_reg[14]) );
  QDFFS gray_avg_reg_reg_2__5_ ( .D(n2757), .CK(clk), .Q(gray_avg_reg[13]) );
  QDFFS gray_avg_reg_reg_2__4_ ( .D(n2756), .CK(clk), .Q(gray_avg_reg[12]) );
  QDFFS gray_avg_reg_reg_2__3_ ( .D(n2755), .CK(clk), .Q(gray_avg_reg[11]) );
  QDFFS gray_avg_reg_reg_2__2_ ( .D(n2754), .CK(clk), .Q(gray_avg_reg[10]) );
  QDFFS gray_avg_reg_reg_2__1_ ( .D(n2753), .CK(clk), .Q(gray_avg_reg[9]) );
  QDFFS gray_avg_reg_reg_2__0_ ( .D(n2752), .CK(clk), .Q(gray_avg_reg[8]) );
  QDFFS gray_avg_reg_reg_3__0_ ( .D(n2751), .CK(clk), .Q(gray_avg_reg[0]) );
  QDFFS gray_avg_reg_reg_3__7_ ( .D(n2750), .CK(clk), .Q(gray_avg_reg[7]) );
  QDFFS gray_avg_reg_reg_3__6_ ( .D(n2749), .CK(clk), .Q(gray_avg_reg[6]) );
  QDFFS gray_avg_reg_reg_3__5_ ( .D(n2748), .CK(clk), .Q(gray_avg_reg[5]) );
  QDFFS gray_avg_reg_reg_3__4_ ( .D(n2747), .CK(clk), .Q(gray_avg_reg[4]) );
  QDFFS gray_avg_reg_reg_3__3_ ( .D(n2746), .CK(clk), .Q(gray_avg_reg[3]) );
  QDFFS gray_avg_reg_reg_3__2_ ( .D(n2745), .CK(clk), .Q(gray_avg_reg[2]) );
  QDFFS gray_avg_reg_reg_3__1_ ( .D(n2744), .CK(clk), .Q(gray_avg_reg[1]) );
  QDFFS SRAM_192X32_data_out_reg_reg_9_ ( .D(n2743), .CK(clk), .Q(
        SRAM_192X32_out_decode[9]) );
  QDFFS SRAM_192X32_data_out_reg_reg_8_ ( .D(n2742), .CK(clk), .Q(
        SRAM_192X32_out_decode[8]) );
  QDFFS SRAM_192X32_data_out_reg_reg_7_ ( .D(n2741), .CK(clk), .Q(
        SRAM_192X32_out_decode[7]) );
  QDFFS SRAM_192X32_data_out_reg_reg_6_ ( .D(n2740), .CK(clk), .Q(
        SRAM_192X32_out_decode[6]) );
  QDFFS SRAM_192X32_data_out_reg_reg_5_ ( .D(n2739), .CK(clk), .Q(
        SRAM_192X32_out_decode[5]) );
  QDFFS SRAM_192X32_data_out_reg_reg_4_ ( .D(n2738), .CK(clk), .Q(
        SRAM_192X32_out_decode[4]) );
  QDFFS SRAM_192X32_data_out_reg_reg_31_ ( .D(n2737), .CK(clk), .Q(
        SRAM_192X32_out_decode[31]) );
  QDFFS SRAM_192X32_data_out_reg_reg_30_ ( .D(n2736), .CK(clk), .Q(
        SRAM_192X32_out_decode[30]) );
  QDFFS SRAM_192X32_data_out_reg_reg_3_ ( .D(n2735), .CK(clk), .Q(
        SRAM_192X32_out_decode[3]) );
  QDFFS SRAM_192X32_data_out_reg_reg_29_ ( .D(n2734), .CK(clk), .Q(
        SRAM_192X32_out_decode[29]) );
  QDFFS SRAM_192X32_data_out_reg_reg_28_ ( .D(n2733), .CK(clk), .Q(
        SRAM_192X32_out_decode[28]) );
  QDFFS SRAM_192X32_data_out_reg_reg_27_ ( .D(n2732), .CK(clk), .Q(
        SRAM_192X32_out_decode[27]) );
  QDFFS SRAM_192X32_data_out_reg_reg_26_ ( .D(n2731), .CK(clk), .Q(
        SRAM_192X32_out_decode[26]) );
  QDFFS SRAM_192X32_data_out_reg_reg_25_ ( .D(n2730), .CK(clk), .Q(
        SRAM_192X32_out_decode[25]) );
  QDFFS SRAM_192X32_data_out_reg_reg_24_ ( .D(n2729), .CK(clk), .Q(
        SRAM_192X32_out_decode[24]) );
  QDFFS SRAM_192X32_data_out_reg_reg_23_ ( .D(n2728), .CK(clk), .Q(
        SRAM_192X32_out_decode[23]) );
  QDFFS SRAM_192X32_data_out_reg_reg_22_ ( .D(n2727), .CK(clk), .Q(
        SRAM_192X32_out_decode[22]) );
  QDFFS SRAM_192X32_data_out_reg_reg_21_ ( .D(n2726), .CK(clk), .Q(
        SRAM_192X32_out_decode[21]) );
  QDFFS SRAM_192X32_data_out_reg_reg_20_ ( .D(n2725), .CK(clk), .Q(
        SRAM_192X32_out_decode[20]) );
  QDFFS SRAM_192X32_data_out_reg_reg_2_ ( .D(n2724), .CK(clk), .Q(
        SRAM_192X32_out_decode[2]) );
  QDFFS SRAM_192X32_data_out_reg_reg_19_ ( .D(n2723), .CK(clk), .Q(
        SRAM_192X32_out_decode[19]) );
  QDFFS SRAM_192X32_data_out_reg_reg_18_ ( .D(n2722), .CK(clk), .Q(
        SRAM_192X32_out_decode[18]) );
  QDFFS SRAM_192X32_data_out_reg_reg_17_ ( .D(n2721), .CK(clk), .Q(
        SRAM_192X32_out_decode[17]) );
  QDFFS SRAM_192X32_data_out_reg_reg_16_ ( .D(n2720), .CK(clk), .Q(
        SRAM_192X32_out_decode[16]) );
  QDFFS SRAM_192X32_data_out_reg_reg_15_ ( .D(n2719), .CK(clk), .Q(
        SRAM_192X32_out_decode[15]) );
  QDFFS SRAM_192X32_data_out_reg_reg_14_ ( .D(n2718), .CK(clk), .Q(
        SRAM_192X32_out_decode[14]) );
  QDFFS SRAM_192X32_data_out_reg_reg_13_ ( .D(n2717), .CK(clk), .Q(
        SRAM_192X32_out_decode[13]) );
  QDFFS SRAM_192X32_data_out_reg_reg_12_ ( .D(n2716), .CK(clk), .Q(
        SRAM_192X32_out_decode[12]) );
  QDFFS SRAM_192X32_data_out_reg_reg_11_ ( .D(n2715), .CK(clk), .Q(
        SRAM_192X32_out_decode[11]) );
  QDFFS SRAM_192X32_data_out_reg_reg_10_ ( .D(n2714), .CK(clk), .Q(
        SRAM_192X32_out_decode[10]) );
  QDFFS SRAM_192X32_data_out_reg_reg_1_ ( .D(n2713), .CK(clk), .Q(
        SRAM_192X32_out_decode[1]) );
  QDFFS SRAM_192X32_data_out_reg_reg_0_ ( .D(n2712), .CK(clk), .Q(
        SRAM_192X32_out_decode[0]) );
  QDFFS filter_result_reg_reg_1__3__7_ ( .D(n2711), .CK(clk), .Q(
        filter_result_reg[39]) );
  QDFFS filter_result_reg_reg_2__3__7_ ( .D(n2710), .CK(clk), .Q(
        filter_result_reg[7]) );
  QDFFS filter_result_reg_reg_1__2__7_ ( .D(n2709), .CK(clk), .Q(
        filter_result_reg[47]) );
  QDFFS filter_result_reg_reg_2__2__7_ ( .D(n2708), .CK(clk), .Q(
        filter_result_reg[15]) );
  QDFFS filter_result_reg_reg_1__1__7_ ( .D(n2707), .CK(clk), .Q(
        filter_result_reg[55]) );
  QDFFS filter_result_reg_reg_2__1__7_ ( .D(n2706), .CK(clk), .Q(
        filter_result_reg[23]) );
  QDFFS filter_result_reg_reg_1__0__7_ ( .D(n2705), .CK(clk), .Q(
        filter_result_reg[63]) );
  QDFFS filter_result_reg_reg_2__0__7_ ( .D(n2704), .CK(clk), .Q(
        filter_result_reg[31]) );
  QDFFS SRAM_64X32_data_out_reg_reg_9_ ( .D(n2703), .CK(clk), .Q(
        SRAM_64X32_out_decode[9]) );
  QDFFS SRAM_64X32_data_out_reg_reg_8_ ( .D(n2702), .CK(clk), .Q(
        SRAM_64X32_out_decode[8]) );
  QDFFS SRAM_64X32_data_out_reg_reg_7_ ( .D(n2701), .CK(clk), .Q(
        SRAM_64X32_out_decode[7]) );
  QDFFS SRAM_64X32_data_out_reg_reg_6_ ( .D(n2700), .CK(clk), .Q(
        SRAM_64X32_out_decode[6]) );
  QDFFS SRAM_64X32_data_out_reg_reg_5_ ( .D(n2699), .CK(clk), .Q(
        SRAM_64X32_out_decode[5]) );
  QDFFS SRAM_64X32_data_out_reg_reg_4_ ( .D(n2698), .CK(clk), .Q(
        SRAM_64X32_out_decode[4]) );
  QDFFS SRAM_64X32_data_out_reg_reg_31_ ( .D(n2697), .CK(clk), .Q(
        SRAM_64X32_out_decode[31]) );
  QDFFS SRAM_64X32_data_out_reg_reg_30_ ( .D(n2696), .CK(clk), .Q(
        SRAM_64X32_out_decode[30]) );
  QDFFS SRAM_64X32_data_out_reg_reg_3_ ( .D(n2695), .CK(clk), .Q(
        SRAM_64X32_out_decode[3]) );
  QDFFS SRAM_64X32_data_out_reg_reg_29_ ( .D(n2694), .CK(clk), .Q(
        SRAM_64X32_out_decode[29]) );
  QDFFS SRAM_64X32_data_out_reg_reg_28_ ( .D(n2693), .CK(clk), .Q(
        SRAM_64X32_out_decode[28]) );
  QDFFS SRAM_64X32_data_out_reg_reg_27_ ( .D(n2692), .CK(clk), .Q(
        SRAM_64X32_out_decode[27]) );
  QDFFS SRAM_64X32_data_out_reg_reg_26_ ( .D(n2691), .CK(clk), .Q(
        SRAM_64X32_out_decode[26]) );
  QDFFS SRAM_64X32_data_out_reg_reg_25_ ( .D(n2690), .CK(clk), .Q(
        SRAM_64X32_out_decode[25]) );
  QDFFS SRAM_64X32_data_out_reg_reg_24_ ( .D(n2689), .CK(clk), .Q(
        SRAM_64X32_out_decode[24]) );
  QDFFS SRAM_64X32_data_out_reg_reg_23_ ( .D(n2688), .CK(clk), .Q(
        SRAM_64X32_out_decode[23]) );
  QDFFS SRAM_64X32_data_out_reg_reg_22_ ( .D(n2687), .CK(clk), .Q(
        SRAM_64X32_out_decode[22]) );
  QDFFS SRAM_64X32_data_out_reg_reg_21_ ( .D(n2686), .CK(clk), .Q(
        SRAM_64X32_out_decode[21]) );
  QDFFS SRAM_64X32_data_out_reg_reg_20_ ( .D(n2685), .CK(clk), .Q(
        SRAM_64X32_out_decode[20]) );
  QDFFS SRAM_64X32_data_out_reg_reg_2_ ( .D(n2684), .CK(clk), .Q(
        SRAM_64X32_out_decode[2]) );
  QDFFS SRAM_64X32_data_out_reg_reg_19_ ( .D(n2683), .CK(clk), .Q(
        SRAM_64X32_out_decode[19]) );
  QDFFS SRAM_64X32_data_out_reg_reg_18_ ( .D(n2682), .CK(clk), .Q(
        SRAM_64X32_out_decode[18]) );
  QDFFS SRAM_64X32_data_out_reg_reg_17_ ( .D(n2681), .CK(clk), .Q(
        SRAM_64X32_out_decode[17]) );
  QDFFS SRAM_64X32_data_out_reg_reg_16_ ( .D(n2680), .CK(clk), .Q(
        SRAM_64X32_out_decode[16]) );
  QDFFS SRAM_64X32_data_out_reg_reg_15_ ( .D(n2679), .CK(clk), .Q(
        SRAM_64X32_out_decode[15]) );
  QDFFS SRAM_64X32_data_out_reg_reg_14_ ( .D(n2678), .CK(clk), .Q(
        SRAM_64X32_out_decode[14]) );
  QDFFS filter_result_reg_reg_1__3__6_ ( .D(n2677), .CK(clk), .Q(
        filter_result_reg[38]) );
  QDFFS filter_result_reg_reg_2__3__6_ ( .D(n2676), .CK(clk), .Q(
        filter_result_reg[6]) );
  QDFFS filter_result_reg_reg_1__2__6_ ( .D(n2675), .CK(clk), .Q(
        filter_result_reg[46]) );
  QDFFS filter_result_reg_reg_2__2__6_ ( .D(n2674), .CK(clk), .Q(
        filter_result_reg[14]) );
  QDFFS filter_result_reg_reg_1__1__6_ ( .D(n2673), .CK(clk), .Q(
        filter_result_reg[54]) );
  QDFFS filter_result_reg_reg_2__1__6_ ( .D(n2672), .CK(clk), .Q(
        filter_result_reg[22]) );
  QDFFS filter_result_reg_reg_1__0__6_ ( .D(n2671), .CK(clk), .Q(
        filter_result_reg[62]) );
  QDFFS filter_result_reg_reg_2__0__6_ ( .D(n2670), .CK(clk), .Q(
        filter_result_reg[30]) );
  QDFFS SRAM_64X32_data_out_reg_reg_13_ ( .D(n2669), .CK(clk), .Q(
        SRAM_64X32_out_decode[13]) );
  QDFFS filter_result_reg_reg_1__3__5_ ( .D(n2668), .CK(clk), .Q(
        filter_result_reg[37]) );
  QDFFS filter_result_reg_reg_2__3__5_ ( .D(n2667), .CK(clk), .Q(
        filter_result_reg[5]) );
  QDFFS filter_result_reg_reg_1__2__5_ ( .D(n2666), .CK(clk), .Q(
        filter_result_reg[45]) );
  QDFFS filter_result_reg_reg_2__2__5_ ( .D(n2665), .CK(clk), .Q(
        filter_result_reg[13]) );
  QDFFS filter_result_reg_reg_1__1__5_ ( .D(n2664), .CK(clk), .Q(
        filter_result_reg[53]) );
  QDFFS filter_result_reg_reg_2__1__5_ ( .D(n2663), .CK(clk), .Q(
        filter_result_reg[21]) );
  QDFFS filter_result_reg_reg_1__0__5_ ( .D(n2662), .CK(clk), .Q(
        filter_result_reg[61]) );
  QDFFS filter_result_reg_reg_2__0__5_ ( .D(n2661), .CK(clk), .Q(
        filter_result_reg[29]) );
  QDFFS SRAM_64X32_data_out_reg_reg_12_ ( .D(n2660), .CK(clk), .Q(
        SRAM_64X32_out_decode[12]) );
  QDFFS filter_result_reg_reg_1__3__4_ ( .D(n2659), .CK(clk), .Q(
        filter_result_reg[36]) );
  QDFFS filter_result_reg_reg_2__3__4_ ( .D(n2658), .CK(clk), .Q(
        filter_result_reg[4]) );
  QDFFS filter_result_reg_reg_1__2__4_ ( .D(n2657), .CK(clk), .Q(
        filter_result_reg[44]) );
  QDFFS filter_result_reg_reg_2__2__4_ ( .D(n2656), .CK(clk), .Q(
        filter_result_reg[12]) );
  QDFFS filter_result_reg_reg_1__1__4_ ( .D(n2655), .CK(clk), .Q(
        filter_result_reg[52]) );
  QDFFS filter_result_reg_reg_2__1__4_ ( .D(n2654), .CK(clk), .Q(
        filter_result_reg[20]) );
  QDFFS filter_result_reg_reg_1__0__4_ ( .D(n2653), .CK(clk), .Q(
        filter_result_reg[60]) );
  QDFFS filter_result_reg_reg_2__0__4_ ( .D(n2652), .CK(clk), .Q(
        filter_result_reg[28]) );
  QDFFS SRAM_64X32_data_out_reg_reg_11_ ( .D(n2651), .CK(clk), .Q(
        SRAM_64X32_out_decode[11]) );
  QDFFS filter_result_reg_reg_1__3__3_ ( .D(n2650), .CK(clk), .Q(
        filter_result_reg[35]) );
  QDFFS filter_result_reg_reg_2__3__3_ ( .D(n2649), .CK(clk), .Q(
        filter_result_reg[3]) );
  QDFFS filter_result_reg_reg_1__2__3_ ( .D(n2648), .CK(clk), .Q(
        filter_result_reg[43]) );
  QDFFS filter_result_reg_reg_2__2__3_ ( .D(n2647), .CK(clk), .Q(
        filter_result_reg[11]) );
  QDFFS filter_result_reg_reg_1__1__3_ ( .D(n2646), .CK(clk), .Q(
        filter_result_reg[51]) );
  QDFFS filter_result_reg_reg_2__1__3_ ( .D(n2645), .CK(clk), .Q(
        filter_result_reg[19]) );
  QDFFS filter_result_reg_reg_1__0__3_ ( .D(n2644), .CK(clk), .Q(
        filter_result_reg[59]) );
  QDFFS filter_result_reg_reg_2__0__3_ ( .D(n2643), .CK(clk), .Q(
        filter_result_reg[27]) );
  QDFFS SRAM_64X32_data_out_reg_reg_10_ ( .D(n2642), .CK(clk), .Q(
        SRAM_64X32_out_decode[10]) );
  QDFFS filter_result_reg_reg_1__3__2_ ( .D(n2641), .CK(clk), .Q(
        filter_result_reg[34]) );
  QDFFS filter_result_reg_reg_2__3__2_ ( .D(n2640), .CK(clk), .Q(
        filter_result_reg[2]) );
  QDFFS filter_result_reg_reg_1__2__2_ ( .D(n2639), .CK(clk), .Q(
        filter_result_reg[42]) );
  QDFFS filter_result_reg_reg_2__2__2_ ( .D(n2638), .CK(clk), .Q(
        filter_result_reg[10]) );
  QDFFS filter_result_reg_reg_1__1__2_ ( .D(n2637), .CK(clk), .Q(
        filter_result_reg[50]) );
  QDFFS filter_result_reg_reg_2__1__2_ ( .D(n2636), .CK(clk), .Q(
        filter_result_reg[18]) );
  QDFFS filter_result_reg_reg_1__0__2_ ( .D(n2635), .CK(clk), .Q(
        filter_result_reg[58]) );
  QDFFS filter_result_reg_reg_2__0__2_ ( .D(n2634), .CK(clk), .Q(
        filter_result_reg[26]) );
  QDFFS SRAM_64X32_data_out_reg_reg_1_ ( .D(n2633), .CK(clk), .Q(
        SRAM_64X32_out_decode[1]) );
  QDFFS filter_result_reg_reg_1__3__1_ ( .D(n2632), .CK(clk), .Q(
        filter_result_reg[33]) );
  QDFFS filter_result_reg_reg_2__3__1_ ( .D(n2631), .CK(clk), .Q(
        filter_result_reg[1]) );
  QDFFS filter_result_reg_reg_1__2__1_ ( .D(n2630), .CK(clk), .Q(
        filter_result_reg[41]) );
  QDFFS filter_result_reg_reg_2__2__1_ ( .D(n2629), .CK(clk), .Q(
        filter_result_reg[9]) );
  QDFFS filter_result_reg_reg_1__1__1_ ( .D(n2628), .CK(clk), .Q(
        filter_result_reg[49]) );
  QDFFS filter_result_reg_reg_2__1__1_ ( .D(n2627), .CK(clk), .Q(
        filter_result_reg[17]) );
  QDFFS filter_result_reg_reg_1__0__1_ ( .D(n2626), .CK(clk), .Q(
        filter_result_reg[57]) );
  QDFFS filter_result_reg_reg_2__0__1_ ( .D(n2625), .CK(clk), .Q(
        filter_result_reg[25]) );
  QDFFS SRAM_64X32_data_out_reg_reg_0_ ( .D(n2624), .CK(clk), .Q(
        SRAM_64X32_out_decode[0]) );
  QDFFS filter_result_reg_reg_1__3__0_ ( .D(n2623), .CK(clk), .Q(
        filter_result_reg[32]) );
  QDFFS filter_result_reg_reg_2__3__0_ ( .D(n2622), .CK(clk), .Q(
        filter_result_reg[0]) );
  QDFFS filter_result_reg_reg_1__2__0_ ( .D(n2621), .CK(clk), .Q(
        filter_result_reg[40]) );
  QDFFS filter_result_reg_reg_2__2__0_ ( .D(n2620), .CK(clk), .Q(
        filter_result_reg[8]) );
  QDFFS filter_result_reg_reg_1__1__0_ ( .D(n2619), .CK(clk), .Q(
        filter_result_reg[48]) );
  QDFFS filter_result_reg_reg_2__1__0_ ( .D(n2618), .CK(clk), .Q(
        filter_result_reg[16]) );
  QDFFS filter_result_reg_reg_1__0__0_ ( .D(n2617), .CK(clk), .Q(
        filter_result_reg[56]) );
  QDFFS filter_result_reg_reg_2__0__0_ ( .D(n2616), .CK(clk), .Q(
        filter_result_reg[24]) );
  QDFFRBS avg_temp_reg_9_ ( .D(n2615), .CK(clk), .RB(rst_n), .Q(avg_temp[9])
         );
  QDFFRBS avg_temp_reg_8_ ( .D(n2614), .CK(clk), .RB(n6308), .Q(avg_temp[8])
         );
  QDFFRBS avg_temp_reg_7_ ( .D(n2613), .CK(clk), .RB(n6308), .Q(avg_temp[7])
         );
  QDFFRBS avg_temp_reg_6_ ( .D(n2612), .CK(clk), .RB(n6307), .Q(avg_temp[6])
         );
  QDFFRBS avg_temp_reg_5_ ( .D(n2611), .CK(clk), .RB(n6308), .Q(avg_temp[5])
         );
  QDFFRBS avg_temp_reg_4_ ( .D(n2610), .CK(clk), .RB(n6308), .Q(avg_temp[4])
         );
  QDFFRBS avg_temp_reg_3_ ( .D(n2609), .CK(clk), .RB(n6308), .Q(avg_temp[3])
         );
  QDFFRBS avg_temp_reg_2_ ( .D(n2608), .CK(clk), .RB(n6306), .Q(avg_temp[2])
         );
  QDFFRBS avg_temp_reg_1_ ( .D(n2607), .CK(clk), .RB(n6307), .Q(avg_temp[1])
         );
  QDFFRBS avg_temp_reg_0_ ( .D(n2606), .CK(clk), .RB(n6308), .Q(avg_temp[0])
         );
  QDFFRBS rd_addr_reg_7_ ( .D(n2605), .CK(clk), .RB(rst_n), .Q(rd_addr[7]) );
  QDFFRBS rd_addr_reg_6_ ( .D(n2604), .CK(clk), .RB(n6308), .Q(rd_addr[6]) );
  QDFFRBS rd_addr_reg_5_ ( .D(n2603), .CK(clk), .RB(n6308), .Q(N1048) );
  QDFFRBS rd_addr_reg_4_ ( .D(n2602), .CK(clk), .RB(n6308), .Q(N1047) );
  QDFFRBS rd_addr_reg_3_ ( .D(n2601), .CK(clk), .RB(n6308), .Q(N1046) );
  QDFFRBS rd_addr_reg_2_ ( .D(n2600), .CK(clk), .RB(n6308), .Q(N1045) );
  QDFFRBS rd_addr_reg_1_ ( .D(n2599), .CK(clk), .RB(n6308), .Q(N1044) );
  QDFFRBS rd_addr_reg_0_ ( .D(n2598), .CK(clk), .RB(n6308), .Q(N1043) );
  QDFFRBS SRAM_192X32_addr_reg_7_ ( .D(n2597), .CK(clk), .RB(rst_n), .Q(
        SRAM_192X32_addr[7]) );
  QDFFRBS SRAM_64X32_addr_reg_0_ ( .D(n2596), .CK(clk), .RB(n6308), .Q(
        SRAM_64X32_addr[0]) );
  QDFFRBS SRAM_64X32_addr_reg_1_ ( .D(n2595), .CK(clk), .RB(n6308), .Q(
        SRAM_64X32_addr[1]) );
  QDFFRBS SRAM_64X32_addr_reg_2_ ( .D(n2594), .CK(clk), .RB(n6308), .Q(
        SRAM_64X32_addr[2]) );
  QDFFRBS SRAM_64X32_addr_reg_3_ ( .D(n2593), .CK(clk), .RB(n6308), .Q(
        SRAM_64X32_addr[3]) );
  QDFFRBS SRAM_64X32_addr_reg_4_ ( .D(n2592), .CK(clk), .RB(n6308), .Q(
        SRAM_64X32_addr[4]) );
  QDFFRBS SRAM_64X32_addr_reg_5_ ( .D(n2591), .CK(clk), .RB(n6308), .Q(
        SRAM_64X32_addr[5]) );
  DFFSBN SRAM_192X32_addr_reg_6_ ( .D(n3206), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[6]), .QB(n6303) );
  DFFSBN wait_conv_out_count_reg_0_ ( .D(n3365), .CK(clk), .SB(n3487), .Q(
        wait_conv_out_count[0]), .QB(n6302) );
  DFFSBN wait_conv_out_count_reg_2_ ( .D(n3364), .CK(clk), .SB(n3487), .Q(
        N6291), .QB(n6304) );
  DFFSBN SRAM_192X32_addr_reg_0_ ( .D(n3212), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[0]) );
  DFFSBN SRAM_192X32_addr_reg_1_ ( .D(n3211), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[1]) );
  DFFSBN SRAM_192X32_addr_reg_2_ ( .D(n3210), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[2]) );
  DFFSBN SRAM_192X32_addr_reg_3_ ( .D(n3209), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[3]) );
  DFFSBN SRAM_192X32_addr_reg_4_ ( .D(n3208), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[4]) );
  DFFSBN SRAM_192X32_addr_reg_5_ ( .D(n3207), .CK(clk), .SB(n3487), .Q(
        SRAM_192X32_addr[5]) );
  QDFFRBN cal_count_reg_2_ ( .D(n3222), .CK(clk), .RB(n6307), .Q(cal_count[2])
         );
  QDFFRBS current_action_idx_reg_0_ ( .D(n3232), .CK(clk), .RB(n6307), .Q(
        current_action_idx[0]) );
  QDFFRBS neg_flag_reg ( .D(n3228), .CK(clk), .RB(n6307), .Q(neg_flag) );
  QDFFRBS find_median_inst_min2_reg_reg_1_ ( .D(find_median_inst_min2[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min2_reg[1]) );
  QDFFRBN find_median_inst_min1_reg_reg_1_ ( .D(find_median_inst_min1[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min1_reg[1]) );
  QDFFRBP wait_conv_out_count_reg_1_ ( .D(n3367), .CK(clk), .RB(n6307), .Q(
        wait_conv_out_count[1]) );
  QDFFRBN find_median_inst_min1_reg_reg_0_ ( .D(find_median_inst_min1[0]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_min1_reg[0]) );
  QDFFRBN out_value_reg ( .D(n2864), .CK(clk), .RB(rst_n), .Q(out_value) );
  QDFFRBN out_valid_reg ( .D(n3196), .CK(clk), .RB(rst_n), .Q(out_valid) );
  QDFFP product_reg_15_ ( .D(N6130), .CK(clk), .Q(product[15]) );
  QDFFRBN flip_flag_reg ( .D(n3371), .CK(clk), .RB(n6306), .Q(flip_flag) );
  QDFFRBN conv_temp_reg_0_ ( .D(n2883), .CK(clk), .RB(rst_n), .Q(conv_temp[0])
         );
  QDFFRBN current_action_idx_reg_1_ ( .D(n3231), .CK(clk), .RB(n6307), .Q(
        current_action_idx[1]) );
  DFFS window_reg_2__2__3_ ( .D(n2965), .CK(clk), .Q(median_in[3]), .QB(n6316)
         );
  DFFS window_reg_2__2__6_ ( .D(n2929), .CK(clk), .Q(median_in[6]), .QB(n6322)
         );
  DFFS image_size_temp_reg_1_ ( .D(n3226), .CK(clk), .Q(image_size_temp[1]), 
        .QB(n3505) );
  QDFFRBN state_reg_0_ ( .D(n3402), .CK(clk), .RB(n6307), .Q(state[0]) );
  QDFFRBN state_reg_3_ ( .D(n3401), .CK(clk), .RB(n6306), .Q(state[3]) );
  QDFFRBS cal_count_reg_7_ ( .D(n3234), .CK(clk), .RB(n6307), .Q(cal_count[7])
         );
  QDFFRBS current_action_idx_reg_2_ ( .D(n3230), .CK(clk), .RB(n6307), .Q(
        current_action_idx[2]) );
  QDFFRBS find_median_inst_max1_reg_reg_1_ ( .D(find_median_inst_max1[1]), 
        .CK(clk), .RB(n6308), .Q(find_median_inst_max1_reg[1]) );
  QDFFRBS cal_count_reg_3_ ( .D(n3223), .CK(clk), .RB(n6307), .Q(cal_count[3])
         );
  QDFFRBS cal_count_reg_1_ ( .D(n3221), .CK(clk), .RB(n6307), .Q(cal_count[1])
         );
  QDFFRBS state_reg_2_ ( .D(n3405), .CK(clk), .RB(n6307), .Q(state[2]) );
  DFFS window_reg_2__2__2_ ( .D(n2977), .CK(clk), .Q(median_in[2]), .QB(n6315)
         );
  DFFS window_reg_2__2__4_ ( .D(n2953), .CK(clk), .Q(median_in[4]), .QB(n6317)
         );
  DFFS window_reg_1__2__2_ ( .D(n2984), .CK(clk), .Q(median_in[26]), .QB(n6318) );
  DFFS window_reg_1__2__1_ ( .D(n2996), .CK(clk), .Q(median_in[25]), .QB(n6310) );
  DFFS window_reg_1__2__6_ ( .D(n2936), .CK(clk), .Q(median_in[30]), .QB(n6312) );
  DFFS window_reg_1__2__4_ ( .D(n2960), .CK(clk), .Q(median_in[28]), .QB(n6311) );
  DFFS window_reg_1__2__3_ ( .D(n2972), .CK(clk), .Q(median_in[27]), .QB(n6319) );
  DFFS window_reg_1__0__2_ ( .D(n2982), .CK(clk), .Q(median_in[42]), .QB(n6313) );
  DFFS window_reg_0__2__5_ ( .D(n2945), .CK(clk), .Q(median_in[53]), .QB(n6321) );
  DFFS window_reg_0__2__0_ ( .D(n3005), .CK(clk), .Q(median_in[48]), .QB(n6320) );
  DFFS window_reg_2__2__1_ ( .D(n2989), .CK(clk), .Q(median_in[1]), .QB(n6314)
         );
  QDFFRBN cal_count_reg_6_ ( .D(n3233), .CK(clk), .RB(n6307), .Q(cal_count[6])
         );
  DFFN image_size_temp_reg_0_ ( .D(n3227), .CK(clk), .Q(image_size_temp[0]), 
        .QB(n6309) );
  QDFFRBN conv_sram_stop_flag_reg_reg ( .D(n6301), .CK(clk), .RB(n6307), .Q(
        conv_sram_stop_flag_reg) );
  INV2 U3574 ( .I(n3889), .O(n4928) );
  MOAI1 U3575 ( .A1(n4304), .A2(n4303), .B1(n5223), .B2(median_in[23]), .O(
        n4312) );
  INV1S U3576 ( .I(n4781), .O(n4921) );
  NR2 U3577 ( .I1(n6190), .I2(n3492), .O(n3899) );
  MAOI1H U3578 ( .A1(n3888), .A2(conv_temp[19]), .B1(n3888), .B2(conv_temp[19]), .O(n3889) );
  INV3 U3579 ( .I(n5520), .O(n5546) );
  MOAI1 U3580 ( .A1(n3835), .A2(n3834), .B1(n3906), .B2(n3907), .O(n3959) );
  BUF2 U3581 ( .I(n4027), .O(n5003) );
  INV3 U3582 ( .I(n5187), .O(n5208) );
  OR2P U3583 ( .I1(n3539), .I2(n3638), .O(n3628) );
  BUF2 U3584 ( .I(n4203), .O(n3485) );
  NR2 U3585 ( .I1(n4542), .I2(SRAM_192_32_read_done), .O(n4081) );
  INV3 U3586 ( .I(n4082), .O(n4542) );
  ND2 U3587 ( .I1(n4945), .I2(n4969), .O(n5745) );
  INV1S U3588 ( .I(state[0]), .O(n5669) );
  INV1S U3589 ( .I(n5746), .O(n5727) );
  INV1S U3590 ( .I(n4119), .O(n3887) );
  INV1S U3591 ( .I(n4580), .O(n4543) );
  ND3S U3592 ( .I1(n3995), .I2(n5755), .I3(n4542), .O(n4034) );
  INV1S U3593 ( .I(state[3]), .O(n4069) );
  INV1S U3594 ( .I(n5753), .O(n3486) );
  ND3S U3595 ( .I1(n4688), .I2(n4432), .I3(n4773), .O(n4981) );
  MOAI1S U3596 ( .A1(n4101), .A2(n4857), .B1(n4095), .B2(n4375), .O(n4698) );
  INV1S U3597 ( .I(n5767), .O(n6245) );
  INV1S U3598 ( .I(n5964), .O(n6032) );
  ND3S U3599 ( .I1(template_count[2]), .I2(n5103), .I3(n5627), .O(n5641) );
  INV1S U3600 ( .I(n3488), .O(n3489) );
  INV1S U3601 ( .I(cal_count[6]), .O(n3488) );
  NR2P U3602 ( .I1(n3492), .I2(n5650), .O(n6196) );
  ND2P U3603 ( .I1(n6003), .I2(n6002), .O(n6004) );
  AO12S U3604 ( .B1(cal_count_5[0]), .B2(n5789), .A1(n5788), .O(n5817) );
  FA1S U3605 ( .A(n5003), .B(N1043), .CI(n4356), .CO(n4368), .S(n4357) );
  AN2 U3606 ( .I1(n5098), .I2(n3666), .O(n5092) );
  XOR2HS U3607 ( .I1(n4031), .I2(n5003), .O(n4356) );
  NR2 U3608 ( .I1(n3902), .I2(n3903), .O(n3881) );
  MAO222 U3609 ( .A1(find_median_inst_min3_reg[7]), .B1(n4355), .C1(n4353), 
        .O(n5397) );
  BUF1 U3610 ( .I(n4448), .O(n4771) );
  ND2 U3611 ( .I1(n6301), .I2(n5712), .O(n5709) );
  ND2 U3612 ( .I1(n5769), .I2(n4512), .O(n4935) );
  ND2 U3613 ( .I1(n5942), .I2(n4105), .O(n4773) );
  BUF1 U3614 ( .I(n4698), .O(n4708) );
  BUF1 U3615 ( .I(n6266), .O(n6263) );
  ND2 U3616 ( .I1(n5727), .I2(n5730), .O(n5738) );
  ND2 U3617 ( .I1(n5728), .I2(n5730), .O(n5739) );
  ND2 U3618 ( .I1(n5729), .I2(n5730), .O(n5740) );
  ND2 U3619 ( .I1(n6243), .I2(n5730), .O(n5742) );
  INV1 U3620 ( .I(n5805), .O(n5860) );
  ND2P U3621 ( .I1(n4386), .I2(n4192), .O(n5934) );
  MOAI1 U3622 ( .A1(n5675), .A2(n4465), .B1(n5675), .B2(n4465), .O(n5861) );
  BUF1 U3623 ( .I(n4647), .O(n5935) );
  ND2 U3624 ( .I1(n4858), .I2(n4857), .O(n5939) );
  MAO222 U3625 ( .A1(n5292), .B1(find_median_inst_max2_reg[7]), .C1(n5291), 
        .O(n5293) );
  MAO222S U3626 ( .A1(n5923), .B1(median_in[30]), .C1(n5140), .O(n5141) );
  NR2P U3627 ( .I1(n5743), .I2(n3647), .O(n6055) );
  INV2 U3628 ( .I(n5259), .O(n5233) );
  MAO222S U3629 ( .A1(n5910), .B1(median_in[29]), .C1(n5139), .O(n5140) );
  ND3 U3630 ( .I1(n3885), .I2(n5918), .I3(n3884), .O(n4782) );
  AN2 U3631 ( .I1(n5591), .I2(n3517), .O(n4956) );
  ND2 U3632 ( .I1(n5635), .I2(n5103), .O(n5637) );
  BUF1 U3633 ( .I(n4786), .O(n4799) );
  INV2 U3634 ( .I(n4788), .O(n4849) );
  INV2 U3635 ( .I(n6210), .O(n6219) );
  MOAI1 U3636 ( .A1(n3887), .A2(n3886), .B1(conv_temp[2]), .B2(product[2]), 
        .O(n4123) );
  ND2 U3637 ( .I1(n5629), .I2(n5101), .O(n5642) );
  ND3 U3638 ( .I1(n5104), .I2(template_count[2]), .I3(n5627), .O(n5639) );
  OR2 U3639 ( .I1(n3676), .I2(n3492), .O(n5626) );
  ND2 U3640 ( .I1(n5636), .I2(n5101), .O(n5644) );
  ND3 U3641 ( .I1(n5636), .I2(template_count[2]), .I3(n5627), .O(n5640) );
  NR2P U3642 ( .I1(n4787), .I2(n5134), .O(n4854) );
  NR2P U3643 ( .I1(n4787), .I2(n5650), .O(n4836) );
  ND2 U3644 ( .I1(n5103), .I2(n5101), .O(n61240) );
  ND2 U3645 ( .I1(n5104), .I2(n5101), .O(n5643) );
  OR2P U3646 ( .I1(n5669), .I2(n5559), .O(n5095) );
  ND2 U3647 ( .I1(n5690), .I2(cal_count[0]), .O(n4608) );
  ND2 U3648 ( .I1(RGB_count[1]), .I2(n3898), .O(n5650) );
  ND3 U3649 ( .I1(n3493), .I2(template_count[3]), .I3(n5102), .O(n5633) );
  AN2 U3650 ( .I1(n5102), .I2(n5627), .O(n5101) );
  OR2S U3651 ( .I1(max_temp[5]), .I2(n5606), .O(n3895) );
  OR2 U3652 ( .I1(RGB_count[1]), .I2(RGB_count[0]), .O(n5610) );
  HA1 U3653 ( .A(product[0]), .B(conv_temp[0]), .C(n4117), .S(n4125) );
  INV1 U3654 ( .I(cal_count[3]), .O(n4945) );
  ND2 U3655 ( .I1(n3505), .I2(n6309), .O(n4553) );
  ND2 U3656 ( .I1(image_size_temp[1]), .I2(image_size_temp[0]), .O(n6242) );
  BUF1 U3657 ( .I(conv_sram_stop_flag_reg), .O(n6265) );
  BUF2 U3658 ( .I(n6308), .O(n3487) );
  INV2 U3659 ( .I(in_valid), .O(n3492) );
  ND2 U3660 ( .I1(n3899), .I2(n5650), .O(n5608) );
  FA1 U3661 ( .A(product[8]), .B(conv_temp[8]), .CI(n4162), .CO(n4164), .S(
        n4163) );
  MOAI1 U3662 ( .A1(n6196), .A2(n6160), .B1(n6196), .B2(n6146), .O(n2839) );
  HA1P U3663 ( .A(image[1]), .B(wgt_temp[0]), .C(n5612), .S(n5611) );
  AOI22H U3664 ( .A1(n5275), .A2(median_in[15]), .B1(n5232), .B2(n4267), .O(
        n5259) );
  NR2T U3665 ( .I1(n5751), .I2(n4627), .O(n4620) );
  INV2 U3666 ( .I(n4746), .O(n5675) );
  ND2 U3667 ( .I1(n5727), .I2(n3547), .O(n3982) );
  INV1CK U3668 ( .I(n3803), .O(n3789) );
  FA1 U3669 ( .A(N1046), .B(n5003), .CI(n4995), .CO(n4992), .S(n4996) );
  FA1 U3670 ( .A(N1047), .B(n5003), .CI(n4992), .CO(n4990), .S(n4993) );
  MOAI1 U3671 ( .A1(n3678), .A2(n3677), .B1(wgt_temp[7]), .B2(n5626), .O(n3354) );
  OAI22H U3672 ( .A1(n4945), .A2(n3983), .B1(n3982), .B2(n4045), .O(n5010) );
  ND2P U3673 ( .I1(n5723), .I2(n5766), .O(n4045) );
  NR2P U3674 ( .I1(n5751), .I2(n3549), .O(n3660) );
  FA1 U3675 ( .A(product[11]), .B(conv_temp[11]), .CI(n4207), .CO(n4111), .S(
        n4208) );
  FA1 U3676 ( .A(product[10]), .B(conv_temp[10]), .CI(n4185), .CO(n4207), .S(
        n4186) );
  FA1 U3677 ( .A(product[13]), .B(conv_temp[13]), .CI(n4113), .CO(n4043), .S(
        n4114) );
  FA1 U3678 ( .A(product[12]), .B(conv_temp[12]), .CI(n4111), .CO(n4113), .S(
        n4112) );
  FA1 U3679 ( .A(product[15]), .B(conv_temp[15]), .CI(n4041), .CO(n4454), .S(
        n4042) );
  FA1 U3680 ( .A(product[14]), .B(conv_temp[14]), .CI(n4043), .CO(n4041), .S(
        n4044) );
  FA1 U3681 ( .A(product[1]), .B(conv_temp[1]), .CI(n4117), .CO(n4119), .S(
        n4118) );
  MOAI1 U3682 ( .A1(n3491), .A2(n4921), .B1(n3491), .B2(conv_out_reg[18]), .O(
        n2857) );
  MOAI1 U3683 ( .A1(n4782), .A2(n4921), .B1(n4956), .B2(conv_temp[18]), .O(
        n2865) );
  MOAI1 U3684 ( .A1(n4782), .A2(n4928), .B1(n4956), .B2(conv_temp[19]), .O(
        n2862) );
  FA1 U3685 ( .A(product[3]), .B(conv_temp[3]), .CI(n4123), .CO(n4115), .S(
        n4124) );
  MOAI1 U3686 ( .A1(n3491), .A2(n4928), .B1(n3491), .B2(conv_out_reg[19]), .O(
        n2858) );
  AO12S U3687 ( .B1(N1047), .B2(n3628), .A1(n3598), .O(n5091) );
  ND2S U3688 ( .I1(n6046), .I2(n5950), .O(n5958) );
  MAO222 U3689 ( .A1(n6043), .B1(pool_temp[12]), .C1(n6020), .O(n6021) );
  MAO222 U3690 ( .A1(pool_temp[11]), .B1(n6040), .C1(n6019), .O(n6020) );
  MAO222 U3691 ( .A1(n6037), .B1(pool_temp[10]), .C1(n6018), .O(n6019) );
  ND2S U3692 ( .I1(n3806), .I2(median_in[11]), .O(n3703) );
  AO12S U3693 ( .B1(N1046), .B2(n3628), .A1(n3605), .O(n5045) );
  ND3S U3694 ( .I1(n3604), .I2(n3603), .I3(n3602), .O(n3605) );
  ND2S U3695 ( .I1(median_in[45]), .I2(n5910), .O(n4282) );
  ND2S U3696 ( .I1(n5869), .I2(n5799), .O(n5808) );
  OR2S U3697 ( .I1(n5679), .I2(n3540), .O(n3577) );
  ND2S U3698 ( .I1(n5729), .I2(cal_count[2]), .O(n4012) );
  ND2S U3699 ( .I1(avg_temp[5]), .I2(n6202), .O(n4217) );
  ND2S U3700 ( .I1(n3547), .I2(n5728), .O(n4604) );
  ND3S U3701 ( .I1(n5954), .I2(n5953), .I3(n5952), .O(n5974) );
  ND2S U3702 ( .I1(n6059), .I2(n5969), .O(n5953) );
  ND3S U3703 ( .I1(n6044), .I2(n5958), .I3(n5951), .O(n5952) );
  MAO222S U3704 ( .A1(n6059), .B1(n5969), .C1(n5968), .O(n5973) );
  ND2S U3705 ( .I1(n6049), .I2(n5967), .O(n5968) );
  MAO222 U3706 ( .A1(pool_temp[21]), .B1(n5875), .C1(n5785), .O(n5786) );
  MAO222 U3707 ( .A1(n5872), .B1(pool_temp[20]), .C1(n5784), .O(n5785) );
  MAO222S U3708 ( .A1(pool_temp[19]), .B1(n5869), .C1(n5783), .O(n5784) );
  MAO222 U3709 ( .A1(n5866), .B1(pool_temp[18]), .C1(n5782), .O(n5783) );
  MAO222S U3710 ( .A1(n5814), .B1(n5858), .C1(n5884), .O(n5829) );
  ND3S U3711 ( .I1(n5796), .I2(n5795), .I3(n5794), .O(n5831) );
  ND2S U3712 ( .I1(n5857), .I2(n5850), .O(n5795) );
  ND3S U3713 ( .I1(n5872), .I2(n5802), .I3(n5793), .O(n5794) );
  FA1S U3714 ( .A(n3868), .B(n3867), .CI(n3866), .CO(n3949), .S(n3951) );
  ND2S U3715 ( .I1(wait_conv_out_count[1]), .I2(n6302), .O(n3679) );
  OR2S U3716 ( .I1(n5020), .I2(n5019), .O(n3508) );
  OR2S U3717 ( .I1(n4945), .I2(n4012), .O(n4016) );
  OR2S U3718 ( .I1(n4003), .I2(n4621), .O(n3996) );
  OR2S U3719 ( .I1(n4009), .I2(n5679), .O(n4033) );
  AN2S U3720 ( .I1(n4008), .I2(n4007), .O(n4009) );
  MAO222 U3721 ( .A1(n5290), .B1(find_median_inst_max2_reg[6]), .C1(n5289), 
        .O(n5291) );
  INV1S U3722 ( .I(n5293), .O(n5294) );
  MAO222 U3723 ( .A1(pool_temp[13]), .B1(n6047), .C1(n6009), .O(n6010) );
  MAO222 U3724 ( .A1(n6044), .B1(pool_temp[12]), .C1(n6008), .O(n6009) );
  MAO222 U3725 ( .A1(pool_temp[11]), .B1(n6041), .C1(n6007), .O(n6008) );
  MAO222 U3726 ( .A1(n6038), .B1(pool_temp[10]), .C1(n6006), .O(n6007) );
  MAO222 U3727 ( .A1(pool_temp[29]), .B1(n6047), .C1(n5979), .O(n5980) );
  MAO222 U3728 ( .A1(n6044), .B1(pool_temp[28]), .C1(n5978), .O(n5979) );
  MAO222 U3729 ( .A1(pool_temp[27]), .B1(n6041), .C1(n5977), .O(n5978) );
  MAO222 U3730 ( .A1(n6038), .B1(pool_temp[26]), .C1(n5976), .O(n5977) );
  OR2S U3731 ( .I1(n4553), .I2(n4191), .O(n5756) );
  ND2S U3732 ( .I1(n4087), .I2(n4092), .O(n4623) );
  ND2S U3733 ( .I1(n4087), .I2(n4942), .O(n4191) );
  AN2S U3734 ( .I1(n5994), .I2(n4986), .O(n5985) );
  ND2S U3735 ( .I1(n4102), .I2(n4386), .O(n4857) );
  AO12S U3736 ( .B1(n4394), .B2(n4393), .A1(n6064), .O(n4510) );
  INV1S U3737 ( .I(neg_flag), .O(n4748) );
  BUF2 U3738 ( .I(n3686), .O(n3806) );
  OR2S U3739 ( .I1(n6302), .I2(wait_conv_out_count[1]), .O(n3685) );
  ND3S U3740 ( .I1(n3684), .I2(wait_conv_out_count[0]), .I3(n6107), .O(n3803)
         );
  INV1 U3741 ( .I(cal_count[1]), .O(n5690) );
  AO12S U3742 ( .B1(N1048), .B2(n3628), .A1(n3594), .O(n5032) );
  AO12S U3743 ( .B1(N1045), .B2(n3628), .A1(n3610), .O(n5058) );
  ND2S U3744 ( .I1(n5092), .I2(N1044), .O(n5074) );
  ND2S U3745 ( .I1(n5092), .I2(N1043), .O(n5086) );
  ND2S U3746 ( .I1(n5093), .I2(SRAM_192X32_addr[0]), .O(n5085) );
  AN2S U3747 ( .I1(n5610), .I2(avg_temp[1]), .O(n6295) );
  AN2S U3748 ( .I1(n5610), .I2(avg_temp[4]), .O(n6283) );
  MAO222S U3749 ( .A1(avg_temp[0]), .B1(avg_temp[1]), .C1(n6206), .O(n4873) );
  AN2S U3750 ( .I1(avg_temp[3]), .I2(n4869), .O(n4870) );
  ND2S U3751 ( .I1(n4638), .I2(n4637), .O(n4639) );
  MAO222S U3752 ( .A1(find_median_inst_min1_reg[1]), .B1(
        find_median_inst_min1_reg[0]), .C1(n4333), .O(n4334) );
  ND2S U3753 ( .I1(n6243), .I2(n3557), .O(n3567) );
  MAO222 U3754 ( .A1(n5284), .B1(find_median_inst_max2_reg[3]), .C1(n5283), 
        .O(n5285) );
  MAO222 U3755 ( .A1(n5282), .B1(find_median_inst_max2_reg[2]), .C1(n5281), 
        .O(n5283) );
  ND2S U3756 ( .I1(median_in[21]), .I2(n5922), .O(n4265) );
  ND2S U3757 ( .I1(n5876), .I2(n5792), .O(n5802) );
  AN2S U3758 ( .I1(n3660), .I2(n4534), .O(n3623) );
  ND2S U3759 ( .I1(n4788), .I2(n5095), .O(n3580) );
  MAO222 U3760 ( .A1(n4341), .B1(find_median_inst_min1_reg[5]), .C1(n4340), 
        .O(n4342) );
  MAO222 U3761 ( .A1(n4339), .B1(find_median_inst_min1_reg[4]), .C1(n4338), 
        .O(n4340) );
  MAO222S U3762 ( .A1(n5893), .B1(median_in[67]), .C1(n5478), .O(n5480) );
  MAO222S U3763 ( .A1(n5528), .B1(median_in[66]), .C1(n5477), .O(n5478) );
  MAO222S U3764 ( .A1(median_in[65]), .B1(median_in[64]), .C1(n5526), .O(n5477) );
  MAO222S U3765 ( .A1(n5460), .B1(find_median_inst_mid_mid_reg[3]), .C1(n5399), 
        .O(n5400) );
  MAO222S U3766 ( .A1(n5457), .B1(find_median_inst_mid_mid_reg[2]), .C1(n5398), 
        .O(n5399) );
  MAO222S U3767 ( .A1(find_median_inst_mid_mid_reg[1]), .B1(
        find_median_inst_mid_mid_reg[0]), .C1(n5430), .O(n5398) );
  ND2S U3768 ( .I1(n5830), .I2(n5832), .O(n5834) );
  AN2S U3769 ( .I1(n5729), .I2(n4969), .O(n5722) );
  HA1S U3770 ( .A(n3859), .B(n3858), .C(n3842), .S(n3946) );
  MOAI1S U3771 ( .A1(n5271), .A2(n3768), .B1(n3799), .B2(median_in[6]), .O(
        n3771) );
  MOAI1S U3772 ( .A1(n5926), .A2(n3767), .B1(n3797), .B2(median_in[38]), .O(
        n3772) );
  OA22S U3773 ( .A1(n4023), .A2(n4022), .B1(n4021), .B2(n4020), .O(n4024) );
  AN2S U3774 ( .I1(cal_count[3]), .I2(n5722), .O(n6240) );
  ND2S U3775 ( .I1(n5721), .I2(n5720), .O(n6244) );
  ND2S U3776 ( .I1(n4226), .I2(avg_temp[6]), .O(n3497) );
  ND2S U3777 ( .I1(avg_temp[8]), .I2(n4210), .O(n4212) );
  AN2S U3778 ( .I1(find_median_inst_max3_reg[5]), .I2(n5310), .O(n5299) );
  MAO222 U3779 ( .A1(n5309), .B1(find_median_inst_max3_reg[4]), .C1(n5297), 
        .O(n5298) );
  MAO222 U3780 ( .A1(find_median_inst_max3_reg[3]), .B1(n5308), .C1(n5296), 
        .O(n5297) );
  ND2S U3781 ( .I1(n5364), .I2(n5363), .O(n5366) );
  MAO222S U3782 ( .A1(find_median_inst_mid1_reg[4]), .B1(n5362), .C1(n5361), 
        .O(n5364) );
  MAO222S U3783 ( .A1(n5378), .B1(find_median_inst_mid1_reg[3]), .C1(n5360), 
        .O(n5361) );
  ND2S U3784 ( .I1(median_in[55]), .I2(n5945), .O(n5541) );
  ND3S U3785 ( .I1(n5326), .I2(n5331), .I3(n5338), .O(n5329) );
  ND2S U3786 ( .I1(n5218), .I2(n5217), .O(n5219) );
  ND2S U3787 ( .I1(n5216), .I2(n5215), .O(n5217) );
  ND2S U3788 ( .I1(n5940), .I2(median_in[71]), .O(n5542) );
  ND2S U3789 ( .I1(median_in[55]), .I2(n5944), .O(n5540) );
  AO12S U3790 ( .B1(median_in[32]), .B2(n5144), .A1(n5143), .O(n4279) );
  AO12S U3791 ( .B1(n5170), .B2(n5169), .A1(n5168), .O(n5171) );
  AN2S U3792 ( .I1(n6028), .I2(n6024), .O(n6016) );
  OA12S U3793 ( .B1(n5975), .B2(n5974), .A1(n5973), .O(n6013) );
  OA12S U3794 ( .B1(n5974), .B2(n5970), .A1(n5973), .O(n6027) );
  ND2S U3795 ( .I1(n5971), .I2(n6034), .O(n5965) );
  ND2S U3796 ( .I1(n5767), .I2(n6242), .O(n4929) );
  ND2S U3797 ( .I1(n5942), .I2(n4093), .O(n4512) );
  ND2S U3798 ( .I1(n4383), .I2(n4378), .O(n4389) );
  ND2S U3799 ( .I1(n5781), .I2(n5994), .O(n5790) );
  MAO222 U3800 ( .A1(n5881), .B1(pool_temp[22]), .C1(n5778), .O(n5780) );
  ND2S U3801 ( .I1(n4087), .I2(n6243), .O(n4378) );
  AN2S U3802 ( .I1(n5757), .I2(n5756), .O(n5764) );
  HA1S U3803 ( .A(n3820), .B(n3819), .C(n3778), .S(n3829) );
  HA1S U3804 ( .A(n3794), .B(n3793), .C(n3866), .S(n3812) );
  ND3S U3805 ( .I1(n4001), .I2(n4000), .I3(n3999), .O(n5680) );
  AO12S U3806 ( .B1(N1044), .B2(n3628), .A1(n3620), .O(n5071) );
  ND2S U3807 ( .I1(n5024), .I2(action_reg_0__0_), .O(n5025) );
  ND3S U3808 ( .I1(n4538), .I2(n4575), .I3(n4537), .O(n4544) );
  ND2S U3809 ( .I1(n4615), .I2(n4614), .O(n5124) );
  ND3S U3810 ( .I1(n4595), .I2(n4594), .I3(n4593), .O(n5131) );
  ND2S U3811 ( .I1(n4630), .I2(n5985), .O(n4593) );
  ND3S U3812 ( .I1(n4590), .I2(n4589), .I3(n4588), .O(n4591) );
  ND3S U3813 ( .I1(n4633), .I2(n4632), .I3(n4631), .O(n5123) );
  ND2S U3814 ( .I1(n5984), .I2(n4630), .O(n4631) );
  ND2S U3815 ( .I1(n5124), .I2(N1043), .O(n5128) );
  AO12S U3816 ( .B1(n3667), .B2(n3628), .A1(n3542), .O(n3585) );
  AO222S U3817 ( .A1(n5727), .A2(n3665), .B1(n5728), .B2(n3664), .C1(n6015), 
        .C2(n3663), .O(n3666) );
  AN2S U3818 ( .I1(n4597), .I2(n3656), .O(n3653) );
  OR3S U3819 ( .I1(n5701), .I2(cal_count_10[3]), .I3(n4033), .O(n4014) );
  AN2S U3820 ( .I1(n5610), .I2(avg_temp[2]), .O(n62910) );
  AN2S U3821 ( .I1(n5610), .I2(avg_temp[5]), .O(n6279) );
  OR2S U3822 ( .I1(n6293), .I2(n6203), .O(n3498) );
  OA12S U3823 ( .B1(avg_temp[4]), .B2(n4224), .A1(n4223), .O(n4871) );
  OAI22S U3824 ( .A1(n5496), .A2(n4320), .B1(n5945), .B2(median_in[63]), .O(
        n5520) );
  MOAI1S U3825 ( .A1(n4319), .A2(n5495), .B1(n4318), .B2(n5490), .O(n4320) );
  ND3S U3826 ( .I1(n4313), .I2(n5485), .I3(n5491), .O(n4317) );
  AN2S U3827 ( .I1(n5994), .I2(cal_count_5[0]), .O(n5984) );
  ND2S U3828 ( .I1(n5013), .I2(n4168), .O(n5712) );
  ND2S U3829 ( .I1(action_idx[1]), .I2(n3991), .O(n4180) );
  AN2S U3830 ( .I1(n4914), .I2(SRAM_out_buffer[56]), .O(n4917) );
  ND2S U3831 ( .I1(n4464), .I2(n4463), .O(n4465) );
  ND2S U3832 ( .I1(n4767), .I2(SRAM_out_buffer[57]), .O(n4975) );
  ND2S U3833 ( .I1(n4767), .I2(SRAM_out_buffer[58]), .O(n4442) );
  ND2S U3834 ( .I1(n4260), .I2(n4259), .O(n4261) );
  ND2S U3835 ( .I1(n4236), .I2(n4235), .O(n4237) );
  OA222S U3836 ( .A1(n5898), .A2(n4894), .B1(n4893), .B2(n5897), .C1(n6041), 
        .C2(n4892), .O(n4980) );
  ND2S U3837 ( .I1(n4233), .I2(n4232), .O(n4234) );
  ND2S U3838 ( .I1(n4767), .I2(SRAM_out_buffer[60]), .O(n5907) );
  ND2S U3839 ( .I1(n4483), .I2(n4482), .O(n4484) );
  ND2S U3840 ( .I1(n4767), .I2(SRAM_out_buffer[61]), .O(n5920) );
  ND2S U3841 ( .I1(n4745), .I2(n4744), .O(n4747) );
  AN2S U3842 ( .I1(n4914), .I2(SRAM_out_buffer[61]), .O(n5912) );
  ND2S U3843 ( .I1(n4205), .I2(n4204), .O(n4206) );
  ND2S U3844 ( .I1(n4767), .I2(SRAM_out_buffer[62]), .O(n4438) );
  AN2S U3845 ( .I1(n4914), .I2(SRAM_out_buffer[62]), .O(n5925) );
  ND2S U3846 ( .I1(n4458), .I2(n4457), .O(n4459) );
  ND2S U3847 ( .I1(n4239), .I2(n4238), .O(n4240) );
  ND2S U3848 ( .I1(n4767), .I2(SRAM_out_buffer[63]), .O(n6065) );
  ND2S U3849 ( .I1(n4254), .I2(n4253), .O(n4255) );
  INV1S U3850 ( .I(n5939), .O(n5943) );
  ND2S U3851 ( .I1(n3537), .I2(state[0]), .O(n3517) );
  AO12S U3852 ( .B1(n5745), .B2(n4466), .A1(n4767), .O(n4504) );
  INV1S U3853 ( .I(n4688), .O(n4772) );
  OR2S U3854 ( .I1(n5770), .I2(n4648), .O(n4416) );
  ND2S U3855 ( .I1(n4257), .I2(n4256), .O(n4258) );
  ND2S U3856 ( .I1(n4248), .I2(n4247), .O(n4249) );
  ND2S U3857 ( .I1(n4421), .I2(n4420), .O(n4422) );
  ND2S U3858 ( .I1(n4245), .I2(n4244), .O(n4246) );
  ND2S U3859 ( .I1(n4425), .I2(n4424), .O(n4426) );
  ND2S U3860 ( .I1(n4251), .I2(n4250), .O(n4252) );
  ND2S U3861 ( .I1(n4451), .I2(n4450), .O(n4452) );
  ND2S U3862 ( .I1(n3806), .I2(median_in[9]), .O(n3687) );
  HA1S U3863 ( .A(n3822), .B(n3821), .C(n3816), .S(n3967) );
  ND3S U3864 ( .I1(n4646), .I2(n4645), .I3(n4644), .O(n2965) );
  ND3S U3865 ( .I1(n4526), .I2(n4525), .I3(n4524), .O(n2989) );
  ND2S U3866 ( .I1(n4889), .I2(window_2__3__1_), .O(n4524) );
  ND3S U3867 ( .I1(n4651), .I2(n4650), .I3(n4649), .O(n2972) );
  ND3S U3868 ( .I1(n4654), .I2(n4653), .I3(n4652), .O(n2960) );
  ND3S U3869 ( .I1(n4657), .I2(n4656), .I3(n4655), .O(n2936) );
  ND3S U3870 ( .I1(n4701), .I2(n4700), .I3(n4699), .O(n2996) );
  ND3S U3871 ( .I1(n4697), .I2(n4696), .I3(n4695), .O(n2984) );
  ND3S U3872 ( .I1(n4694), .I2(n4693), .I3(n4692), .O(n2953) );
  AO22S U3873 ( .A1(n3493), .A2(n6296), .B1(n3492), .B2(avg_temp[1]), .O(n2607) );
  MAO222 U3874 ( .A1(find_median_inst_max2_reg[1]), .B1(
        find_median_inst_max2_reg[0]), .C1(n5280), .O(n5281) );
  MAO222 U3875 ( .A1(n4337), .B1(find_median_inst_min1_reg[3]), .C1(n4336), 
        .O(n4338) );
  MAO222 U3876 ( .A1(n4335), .B1(find_median_inst_min1_reg[2]), .C1(n4334), 
        .O(n4336) );
  AO22S U3877 ( .A1(pool_temp[2]), .A2(n5866), .B1(n5835), .B2(n3513), .O(
        n3514) );
  OR2S U3878 ( .I1(pool_temp[2]), .I2(n5866), .O(n3513) );
  MAO222 U3879 ( .A1(n5860), .B1(n5863), .C1(pool_temp[1]), .O(n5835) );
  MAO222 U3880 ( .A1(n5860), .B1(n5863), .C1(pool_temp[17]), .O(n5782) );
  OR2S U3881 ( .I1(n5746), .I2(n4103), .O(n5749) );
  ND2S U3882 ( .I1(n3568), .I2(n3558), .O(n4585) );
  OR2S U3883 ( .I1(n3570), .I2(n3569), .O(n4532) );
  ND2S U3884 ( .I1(n4625), .I2(n4528), .O(n4602) );
  OR2S U3885 ( .I1(n3570), .I2(n5758), .O(n4555) );
  OR2S U3886 ( .I1(n4582), .I2(n4562), .O(n4552) );
  AN2S U3887 ( .I1(n4620), .I2(n4534), .O(n4587) );
  ND2S U3888 ( .I1(n4546), .I2(n4545), .O(n4548) );
  OR2S U3889 ( .I1(n4530), .I2(n5679), .O(n4531) );
  AN2S U3890 ( .I1(n3657), .I2(n4545), .O(n3561) );
  NR2 U3891 ( .I1(n6299), .I2(n5654), .O(n3657) );
  ND2 U3892 ( .I1(n3537), .I2(n3657), .O(n3549) );
  ND2 U3893 ( .I1(n4358), .I2(n5678), .O(n4547) );
  INV1S U3894 ( .I(n4094), .O(n4002) );
  MAO222S U3895 ( .A1(n5602), .B1(max_temp[1]), .C1(n5601), .O(n3890) );
  ND2S U3896 ( .I1(median_in[69]), .I2(n5914), .O(n4315) );
  MAO222 U3897 ( .A1(n5288), .B1(find_median_inst_max2_reg[5]), .C1(n5287), 
        .O(n5289) );
  MAO222 U3898 ( .A1(n5286), .B1(find_median_inst_max2_reg[4]), .C1(n5285), 
        .O(n5287) );
  MAO222 U3899 ( .A1(n5307), .B1(find_median_inst_max3_reg[2]), .C1(n5295), 
        .O(n5296) );
  MAO222 U3900 ( .A1(n5306), .B1(find_median_inst_max3_reg[1]), .C1(n5305), 
        .O(n5295) );
  MAO222S U3901 ( .A1(n5376), .B1(find_median_inst_mid2_reg[3]), .C1(n5322), 
        .O(n5332) );
  MAO222S U3902 ( .A1(n5373), .B1(find_median_inst_mid2_reg[2]), .C1(n5321), 
        .O(n5322) );
  MAO222S U3903 ( .A1(find_median_inst_mid2_reg[1]), .B1(
        find_median_inst_mid2_reg[0]), .C1(n5320), .O(n5321) );
  ND2S U3904 ( .I1(n5368), .I2(find_median_inst_mid2_reg[7]), .O(n5339) );
  MAO222S U3905 ( .A1(median_in[4]), .B1(n5906), .C1(n5214), .O(n5216) );
  MAO222S U3906 ( .A1(n5267), .B1(median_in[3]), .C1(n5213), .O(n5214) );
  MAO222S U3907 ( .A1(n5265), .B1(median_in[2]), .C1(n5212), .O(n5213) );
  MAO222S U3908 ( .A1(median_in[1]), .B1(median_in[0]), .C1(n5263), .O(n5212)
         );
  ND2S U3909 ( .I1(n4263), .I2(n4265), .O(n5229) );
  MOAI1S U3910 ( .A1(median_in[18]), .A2(n5265), .B1(n5268), .B2(median_in[11]), .O(n5226) );
  MOAI1S U3911 ( .A1(median_in[41]), .A2(n5177), .B1(n6313), .B2(median_in[34]), .O(n5143) );
  OR3S U3912 ( .I1(n4281), .I2(n5185), .I3(median_in[36]), .O(n4280) );
  ND2 U3913 ( .I1(n4004), .I2(n4002), .O(n3984) );
  ND2S U3914 ( .I1(wait_conv_out_count[3]), .I2(N6291), .O(n6083) );
  ND3S U3915 ( .I1(n5959), .I2(n5958), .I3(n5957), .O(n5972) );
  ND2S U3916 ( .I1(n3489), .I2(cal_count[7]), .O(n5750) );
  ND2S U3917 ( .I1(n5745), .I2(n5727), .O(n4096) );
  MAO222 U3918 ( .A1(n5878), .B1(pool_temp[6]), .C1(n5838), .O(n5839) );
  MAO222S U3919 ( .A1(pool_temp[5]), .B1(n5875), .C1(n5837), .O(n5838) );
  MAO222 U3920 ( .A1(n5872), .B1(pool_temp[4]), .C1(n5836), .O(n5837) );
  MAO222 U3921 ( .A1(pool_temp[3]), .B1(n5869), .C1(n3514), .O(n5836) );
  MAO222 U3922 ( .A1(pool_temp[21]), .B1(n5876), .C1(n5777), .O(n5778) );
  MAO222 U3923 ( .A1(pool_temp[20]), .B1(n5873), .C1(n5776), .O(n5777) );
  MAO222 U3924 ( .A1(n5870), .B1(pool_temp[19]), .C1(n5775), .O(n5776) );
  MAO222 U3925 ( .A1(pool_temp[18]), .B1(n5867), .C1(n5774), .O(n5775) );
  ND2S U3926 ( .I1(n5809), .I2(n5808), .O(n5830) );
  ND3S U3927 ( .I1(n5867), .I2(n5808), .I3(n5800), .O(n5801) );
  ND2S U3928 ( .I1(n4509), .I2(n4379), .O(n4393) );
  ND2S U3929 ( .I1(n4102), .I2(n4101), .O(n4394) );
  ND3S U3930 ( .I1(n6093), .I2(n3684), .I3(n6302), .O(n3769) );
  OR2S U3931 ( .I1(n6071), .I2(n6114), .O(n3768) );
  ND2S U3932 ( .I1(n3806), .I2(median_in[12]), .O(n3726) );
  AN2S U3933 ( .I1(n6243), .I2(n4376), .O(n4092) );
  ND2 U3934 ( .I1(n5669), .I2(n5010), .O(n3992) );
  ND2S U3935 ( .I1(n5766), .I2(n5680), .O(n4056) );
  AO12S U3936 ( .B1(N1048), .B2(n3641), .A1(n3595), .O(n3596) );
  AO12S U3937 ( .B1(n3639), .B2(SRAM_192X32_addr[5]), .A1(n3637), .O(n3595) );
  AO12S U3938 ( .B1(N1047), .B2(n3641), .A1(n3599), .O(n3600) );
  AO12S U3939 ( .B1(n3639), .B2(SRAM_192X32_addr[4]), .A1(n3637), .O(n3599) );
  AO12S U3940 ( .B1(N1046), .B2(n3641), .A1(n3606), .O(n3607) );
  AO12S U3941 ( .B1(n3639), .B2(SRAM_192X32_addr[3]), .A1(n3637), .O(n3606) );
  AO12S U3942 ( .B1(N1045), .B2(n3641), .A1(n3611), .O(n3612) );
  AO12S U3943 ( .B1(N1044), .B2(n3641), .A1(n3640), .O(n3642) );
  AO12S U3944 ( .B1(N1043), .B2(n3628), .A1(n3627), .O(n5079) );
  ND2S U3945 ( .I1(n3547), .I2(n3525), .O(n4613) );
  OR2S U3946 ( .I1(n4563), .I2(n4562), .O(n4573) );
  OR2S U3947 ( .I1(n4566), .I2(n4565), .O(n4630) );
  OA12S U3948 ( .B1(n4618), .B2(n4617), .A1(n4616), .O(n4622) );
  AO12S U3949 ( .B1(n5026), .B2(n3641), .A1(n3588), .O(n3589) );
  ND3S U3950 ( .I1(n3587), .I2(n3630), .I3(n3586), .O(n3588) );
  AO12S U3951 ( .B1(n5026), .B2(n3628), .A1(n3592), .O(n5019) );
  AO12S U3952 ( .B1(n3667), .B2(n3641), .A1(n3582), .O(n3583) );
  OR2S U3953 ( .I1(n3486), .I2(n3549), .O(n3662) );
  ND2S U3954 ( .I1(n4025), .I2(n4012), .O(n4554) );
  ND2S U3955 ( .I1(cal_count_5[2]), .I2(n3645), .O(n3646) );
  AN2S U3956 ( .I1(n3995), .I2(n5729), .O(n4019) );
  OR2S U3957 ( .I1(n4621), .I2(n4392), .O(n4025) );
  MAO222 U3958 ( .A1(n5605), .B1(max_temp[4]), .C1(n3894), .O(n3896) );
  MAO222 U3959 ( .A1(n5604), .B1(max_temp[3]), .C1(n3893), .O(n3894) );
  MOAI1S U3960 ( .A1(n3892), .A2(n3891), .B1(max_temp[2]), .B2(n5603), .O(
        n3893) );
  INV1S U3961 ( .I(n3890), .O(n3892) );
  ND2S U3962 ( .I1(median_in[58]), .I2(n5533), .O(n5487) );
  ND2S U3963 ( .I1(median_in[67]), .I2(n5895), .O(n5490) );
  OR3B2S U3964 ( .I1(n4319), .B1(n4316), .B2(n4315), .O(n5492) );
  OR3S U3965 ( .I1(n4314), .I2(n5532), .I3(median_in[60]), .O(n4316) );
  ND2S U3966 ( .I1(median_in[59]), .I2(n5894), .O(n5494) );
  MAO222 U3967 ( .A1(n4345), .B1(find_median_inst_min1_reg[7]), .C1(n4344), 
        .O(n4346) );
  MAO222 U3968 ( .A1(n4343), .B1(find_median_inst_min1_reg[6]), .C1(n4342), 
        .O(n4344) );
  INV1S U3969 ( .I(n4346), .O(n4347) );
  MAO222 U3970 ( .A1(n5393), .B1(find_median_inst_min3_reg[3]), .C1(n4349), 
        .O(n4350) );
  MAO222 U3971 ( .A1(find_median_inst_min3_reg[2]), .B1(n5392), .C1(n4348), 
        .O(n4349) );
  MAO222 U3972 ( .A1(find_median_inst_min3_reg[1]), .B1(n4354), .C1(n5391), 
        .O(n4348) );
  AO12S U3973 ( .B1(n5271), .B2(median_in[6]), .A1(n5255), .O(n5252) );
  AO12S U3974 ( .B1(n5484), .B2(n5483), .A1(n5482), .O(n5502) );
  ND2S U3975 ( .I1(n5481), .I2(n5541), .O(n5482) );
  ND3S U3976 ( .I1(n5439), .I2(n5444), .I3(n5438), .O(n5440) );
  AO12S U3977 ( .B1(n5404), .B2(n5403), .A1(n5402), .O(n5405) );
  HA1 U3978 ( .A(conv_temp[16]), .B(n4454), .C(n4713), .S(n4455) );
  FA1S U3979 ( .A(product[9]), .B(conv_temp[9]), .CI(n4164), .CO(n4185), .S(
        n4165) );
  FA1S U3980 ( .A(product[6]), .B(conv_temp[6]), .CI(n4126), .CO(n4155), .S(
        n4127) );
  FA1S U3981 ( .A(product[5]), .B(conv_temp[5]), .CI(n4121), .CO(n4126), .S(
        n4122) );
  ND2S U3982 ( .I1(cal_count[1]), .I2(n5725), .O(n3516) );
  ND2S U3983 ( .I1(n5744), .I2(n4056), .O(n5678) );
  ND2S U3984 ( .I1(action_idx[2]), .I2(n5579), .O(n5568) );
  ND2S U3985 ( .I1(n61230), .I2(n5572), .O(n5567) );
  ND2S U3986 ( .I1(template_count[0]), .I2(template_count[1]), .O(n5100) );
  ND2S U3987 ( .I1(n5753), .I2(n4088), .O(n4931) );
  AN2S U3988 ( .I1(n4096), .I2(n5755), .O(n4388) );
  MAO222 U3989 ( .A1(n5857), .B1(pool_temp[23]), .C1(n5787), .O(n5789) );
  MAO222 U3990 ( .A1(n5878), .B1(pool_temp[22]), .C1(n5786), .O(n5787) );
  ND2S U3991 ( .I1(n6243), .I2(n4375), .O(n4391) );
  ND2S U3992 ( .I1(n4945), .I2(n5722), .O(n4387) );
  ND2S U3993 ( .I1(n4191), .I2(n5725), .O(n4229) );
  ND2S U3994 ( .I1(n6240), .I2(n5723), .O(n5724) );
  ND2S U3995 ( .I1(n3991), .I2(n5576), .O(n4988) );
  FA1S U3996 ( .A(n3809), .B(n3808), .CI(n3807), .CO(n3872), .S(n3815) );
  FA1S U3997 ( .A(n3946), .B(n3945), .CI(n3944), .CO(n3975), .S(n3978) );
  FA1S U3998 ( .A(n3877), .B(n3876), .CI(n3875), .CO(n3878), .S(n3973) );
  ND2S U3999 ( .I1(n3806), .I2(median_in[14]), .O(n3774) );
  ND3S U4000 ( .I1(n3763), .I2(n3762), .I3(n3761), .O(n3766) );
  AN2S U4001 ( .I1(n5632), .I2(template_count[1]), .O(n5104) );
  AN2S U4002 ( .I1(n5678), .I2(n4076), .O(n4157) );
  INV1S U4003 ( .I(n4608), .O(n5728) );
  AN2S U4004 ( .I1(n6243), .I2(n4003), .O(n4942) );
  ND2S U4005 ( .I1(n4358), .I2(n4157), .O(n4160) );
  OR2S U4006 ( .I1(wait_conv_out_count[0]), .I2(wait_conv_out_count[1]), .O(
        n6071) );
  MOAI1S U4007 ( .A1(n5546), .A2(median_in[57]), .B1(n5546), .B2(n5534), .O(
        n5548) );
  MOAI1S U4008 ( .A1(n5208), .A2(median_in[33]), .B1(n5208), .B2(n5188), .O(
        n5198) );
  INV1S U4009 ( .I(n4090), .O(n4967) );
  ND2S U4010 ( .I1(n5918), .I2(n5558), .O(n4168) );
  FA1S U4011 ( .A(N1045), .B(n4999), .CI(n4998), .CO(n4995), .S(n5000) );
  AO112S U4012 ( .C1(n4037), .C2(n5984), .A1(n4010), .B1(n4013), .O(n4011) );
  FA1S U4013 ( .A(N1048), .B(n5003), .CI(n4990), .CO(n5002), .S(n4039) );
  HA1S U4014 ( .A(image[0]), .B(n6297), .C(n6294), .S(n6298) );
  AN2S U4015 ( .I1(n5610), .I2(avg_temp[0]), .O(n6297) );
  AN2S U4016 ( .I1(n5610), .I2(avg_temp[3]), .O(n6287) );
  AN2S U4017 ( .I1(n5610), .I2(avg_temp[6]), .O(n6275) );
  ND2S U4018 ( .I1(avg_temp[5]), .I2(n4218), .O(n4215) );
  MAO222 U4019 ( .A1(n5609), .B1(max_temp[7]), .C1(n3897), .O(n6190) );
  MAO222 U4020 ( .A1(n3900), .B1(max_temp[6]), .C1(n3490), .O(n3897) );
  AO22S U4021 ( .A1(max_temp[5]), .A2(n5606), .B1(n3896), .B2(n3895), .O(n3490) );
  HA1S U4022 ( .A(image[2]), .B(wgt_temp[0]), .C(n6157), .S(n6159) );
  MOAI1S U4023 ( .A1(n5233), .A2(median_in[9]), .B1(n5233), .B2(n5264), .O(
        n4307) );
  MOAI1S U4024 ( .A1(n5208), .A2(median_in[41]), .B1(n5208), .B2(n5177), .O(
        n4296) );
  ND2S U4025 ( .I1(n5466), .I2(n5468), .O(n5471) );
  MOAI1 U4026 ( .A1(find_median_inst_max3_reg[7]), .A2(n5304), .B1(n5313), 
        .B2(n5303), .O(n5312) );
  MAO222S U4027 ( .A1(find_median_inst_max3_reg[6]), .B1(n5311), .C1(n5302), 
        .O(n5304) );
  AO22 U4028 ( .A1(n6067), .A2(n5255), .B1(n4785), .B2(n4273), .O(n5279) );
  MAO222S U4029 ( .A1(n4276), .B1(median_in[6]), .C1(n4272), .O(n4273) );
  MAO222 U4030 ( .A1(n5278), .B1(median_in[5]), .C1(n4271), .O(n4272) );
  MAO222 U4031 ( .A1(n4277), .B1(median_in[4]), .C1(n4270), .O(n4271) );
  MAO222 U4032 ( .A1(find_median_inst_min3_reg[6]), .B1(n5396), .C1(n4352), 
        .O(n4353) );
  MAO222 U4033 ( .A1(find_median_inst_min3_reg[5]), .B1(n5395), .C1(n4351), 
        .O(n4352) );
  MAO222 U4034 ( .A1(find_median_inst_min3_reg[4]), .B1(n5394), .C1(n4350), 
        .O(n4351) );
  OR2S U4035 ( .I1(n5255), .I2(n5221), .O(n4303) );
  MAO222S U4036 ( .A1(n4306), .B1(median_in[6]), .C1(n4302), .O(n4304) );
  MAO222 U4037 ( .A1(n4311), .B1(median_in[5]), .C1(n4301), .O(n4302) );
  MAO222S U4038 ( .A1(find_median_inst_mid3_reg[7]), .B1(n5368), .C1(n5367), 
        .O(n5370) );
  ND2S U4039 ( .I1(n5382), .I2(n5384), .O(n5387) );
  MOAI1 U4040 ( .A1(median_in[63]), .A2(n5541), .B1(n4784), .B2(n4326), .O(
        n5556) );
  MAO222S U4041 ( .A1(n5555), .B1(median_in[54]), .C1(n4325), .O(n4326) );
  MAO222 U4042 ( .A1(n4328), .B1(median_in[53]), .C1(n4324), .O(n4325) );
  MAO222 U4043 ( .A1(median_in[52]), .B1(n4330), .C1(n4323), .O(n4324) );
  ND2S U4044 ( .I1(n5541), .I2(n5540), .O(n5543) );
  MAO222S U4045 ( .A1(median_in[54]), .B1(n5553), .C1(n5539), .O(n5544) );
  MAO222 U4046 ( .A1(n5552), .B1(median_in[53]), .C1(n5538), .O(n5539) );
  MAO222 U4047 ( .A1(median_in[31]), .B1(n4292), .C1(n4291), .O(n5211) );
  MAO222 U4048 ( .A1(median_in[30]), .B1(n4294), .C1(n4290), .O(n4291) );
  MAO222 U4049 ( .A1(n5210), .B1(median_in[29]), .C1(n4289), .O(n4290) );
  OAI22S U4050 ( .A1(n5936), .A2(n5196), .B1(median_in[31]), .B2(n5195), .O(
        n5204) );
  ND2S U4051 ( .I1(median_in[47]), .I2(n5194), .O(n5196) );
  ND2S U4052 ( .I1(median_in[31]), .I2(n5195), .O(n5194) );
  MAO222S U4053 ( .A1(median_in[30]), .B1(n5203), .C1(n5193), .O(n5195) );
  ND2S U4054 ( .I1(n5369), .I2(n5330), .O(n5356) );
  OR2S U4055 ( .I1(n5223), .I2(n5222), .O(n5234) );
  MAO222S U4056 ( .A1(n5219), .B1(n5270), .C1(median_in[6]), .O(n5220) );
  ND2S U4057 ( .I1(n5272), .I2(n5273), .O(n5274) );
  OA12S U4058 ( .B1(n5519), .B2(n5518), .A1(n5540), .O(n5521) );
  ND2S U4059 ( .I1(n5529), .I2(n5530), .O(n5531) );
  MAO222S U4060 ( .A1(n5936), .B1(median_in[31]), .C1(n5141), .O(n5151) );
  ND2S U4061 ( .I1(n5173), .I2(n5171), .O(n5172) );
  ND2S U4062 ( .I1(median_in[31]), .I2(n5205), .O(n5173) );
  ND2S U4063 ( .I1(n5180), .I2(n5181), .O(n5182) );
  AN2S U4064 ( .I1(find_median_inst_max2_reg[7]), .I2(
        find_median_inst_max1_reg[7]), .O(n5313) );
  ND2S U4065 ( .I1(cal_count_5[2]), .I2(n6028), .O(n5713) );
  ND2S U4066 ( .I1(cal_count_5[0]), .I2(n5714), .O(n5710) );
  AO12S U4067 ( .B1(n4987), .B2(n4986), .A1(n5695), .O(n5711) );
  ND2S U4068 ( .I1(n5697), .I2(n5700), .O(n5702) );
  ND2S U4069 ( .I1(n5707), .I2(n5704), .O(n5697) );
  ND2S U4070 ( .I1(n5715), .I2(n5696), .O(n5704) );
  OR2S U4071 ( .I1(cal_count[4]), .I2(n4942), .O(n5688) );
  ND2S U4072 ( .I1(cal_count[4]), .I2(n4942), .O(n5687) );
  OA12S U4073 ( .B1(n4985), .B2(n5655), .A1(n6301), .O(n5657) );
  ND2S U4074 ( .I1(n5767), .I2(n5010), .O(n5667) );
  FA1S U4075 ( .A(image[4]), .B(wgt_temp[3]), .CI(n5616), .CO(n5618), .S(n5617) );
  FA1S U4076 ( .A(image[2]), .B(wgt_temp[1]), .CI(n5612), .CO(n5614), .S(n5613) );
  INV1S U4077 ( .I(image[1]), .O(n5602) );
  INV1S U4078 ( .I(image[0]), .O(n5601) );
  NR2 U4079 ( .I1(n6196), .I2(n3899), .O(n5607) );
  ND2S U4080 ( .I1(RGB_count[0]), .I2(n3675), .O(n5134) );
  OA12S U4081 ( .B1(n5669), .B2(n5133), .A1(n3492), .O(n5135) );
  ND2S U4082 ( .I1(n4962), .I2(n5593), .O(n4952) );
  AN2S U4083 ( .I1(n5567), .I2(n5568), .O(n5569) );
  ND2S U4084 ( .I1(action_idx[0]), .I2(in_valid2), .O(n5566) );
  ND2S U4085 ( .I1(n5566), .I2(n5567), .O(n5565) );
  OR2S U4086 ( .I1(state[0]), .I2(n5559), .O(n5591) );
  NR2 U4087 ( .I1(template_count[3]), .I2(n3492), .O(n5627) );
  ND2S U4088 ( .I1(SRAM_out_buffer[56]), .I2(n4767), .O(n4983) );
  ND2S U4089 ( .I1(n4690), .I2(n4689), .O(n4691) );
  INV1S U4090 ( .I(median_in[61]), .O(n5914) );
  AOI22S U4091 ( .A1(n6017), .A2(n6016), .B1(n6015), .B2(n6014), .O(n6051) );
  MAO222 U4092 ( .A1(pool_temp[15]), .B1(n6059), .C1(n6011), .O(n6012) );
  MAO222 U4093 ( .A1(n6052), .B1(pool_temp[14]), .C1(n6010), .O(n6011) );
  ND3 U4094 ( .I1(n6028), .I2(n6027), .I3(n6026), .O(n6050) );
  MAO222 U4095 ( .A1(pool_temp[15]), .B1(n6029), .C1(n6023), .O(n6025) );
  MAO222 U4096 ( .A1(n6049), .B1(pool_temp[14]), .C1(n6022), .O(n6023) );
  ND2P U4097 ( .I1(n6051), .I2(n6050), .O(n6053) );
  MAO222 U4098 ( .A1(pool_temp[31]), .B1(n6059), .C1(n5981), .O(n5982) );
  MAO222 U4099 ( .A1(n6052), .B1(pool_temp[30]), .C1(n5980), .O(n5981) );
  MAO222 U4100 ( .A1(n6049), .B1(pool_temp[30]), .C1(n5990), .O(n5991) );
  ND2S U4101 ( .I1(n5856), .I2(n5852), .O(n5882) );
  AOI13HS U4102 ( .B1(n5854), .B2(cal_count_5[2]), .B3(n6028), .A1(n5853), .O(
        n5880) );
  OR2B1S U4103 ( .I1(n5856), .B1(n5855), .O(n5879) );
  ND2S U4104 ( .I1(cal_count_5[2]), .I2(n5854), .O(n5855) );
  OR3B2S U4105 ( .I1(n5770), .B1(n5769), .B2(n5768), .O(n5773) );
  ND2S U4106 ( .I1(n4198), .I2(n4197), .O(n4199) );
  ND2S U4107 ( .I1(n4108), .I2(n4107), .O(n4109) );
  ND2S U4108 ( .I1(n4480), .I2(n4479), .O(n4481) );
  ND2S U4109 ( .I1(n5758), .I2(n5762), .O(n5760) );
  ND2S U4110 ( .I1(n4471), .I2(n4470), .O(n4472) );
  INV1S U4111 ( .I(n6060), .O(n5931) );
  ND2S U4112 ( .I1(n5582), .I2(in_valid2), .O(n5583) );
  OR2S U4113 ( .I1(n4988), .I2(n5572), .O(n4989) );
  OR2S U4114 ( .I1(n5585), .I2(n5584), .O(n5589) );
  ND2S U4115 ( .I1(n5580), .I2(n5579), .O(n5581) );
  OR2S U4116 ( .I1(n5584), .I2(n5574), .O(n5575) );
  ND2S U4117 ( .I1(n5577), .I2(n5576), .O(n5578) );
  ND2S U4118 ( .I1(action_idx[1]), .I2(n5577), .O(n5573) );
  FA1S U4119 ( .A(n3818), .B(n3817), .CI(n3816), .CO(n3833), .S(n3964) );
  FA1S U4120 ( .A(n3830), .B(n3829), .CI(n3828), .CO(n3907), .S(n3963) );
  ND3S U4121 ( .I1(n3788), .I2(n3787), .I3(n3786), .O(n3792) );
  ND3S U4122 ( .I1(n3802), .I2(n3801), .I3(n3800), .O(n3805) );
  ND2S U4123 ( .I1(n5627), .I2(n5631), .O(n5638) );
  ND3S U4124 ( .I1(n4515), .I2(n4514), .I3(n4513), .O(n3005) );
  ND2S U4125 ( .I1(n4889), .I2(window_0__3__0_), .O(n4514) );
  ND2S U4126 ( .I1(n4903), .I2(n4902), .O(n2945) );
  ND2S U4127 ( .I1(n4970), .I2(n3517), .O(n4973) );
  AO12S U4128 ( .B1(n5036), .B2(n5098), .A1(n5035), .O(n3207) );
  ND2S U4129 ( .I1(n5093), .I2(SRAM_192X32_addr[5]), .O(n5033) );
  ND2S U4130 ( .I1(n5092), .I2(N1048), .O(n5034) );
  AO12S U4131 ( .B1(n5099), .B2(n5098), .A1(n5097), .O(n3208) );
  ND2S U4132 ( .I1(n5093), .I2(SRAM_192X32_addr[4]), .O(n5094) );
  ND2S U4133 ( .I1(n5092), .I2(N1047), .O(n5096) );
  AO12S U4134 ( .B1(n5049), .B2(n5098), .A1(n5048), .O(n3209) );
  ND2S U4135 ( .I1(n5093), .I2(SRAM_192X32_addr[3]), .O(n5046) );
  ND2S U4136 ( .I1(n5092), .I2(N1046), .O(n5047) );
  AO12S U4137 ( .B1(n5062), .B2(n5098), .A1(n5061), .O(n3210) );
  ND2S U4138 ( .I1(n5093), .I2(SRAM_192X32_addr[2]), .O(n5059) );
  ND2S U4139 ( .I1(n5092), .I2(N1045), .O(n5060) );
  AO12S U4140 ( .B1(n5076), .B2(n5098), .A1(n5075), .O(n3211) );
  ND2S U4141 ( .I1(n5093), .I2(SRAM_192X32_addr[1]), .O(n5073) );
  AO12S U4142 ( .B1(n5088), .B2(n5098), .A1(n5087), .O(n3212) );
  ND2S U4143 ( .I1(n5092), .I2(n5026), .O(n5027) );
  ND2S U4144 ( .I1(n5123), .I2(wb_addr[5]), .O(n5118) );
  ND2S U4145 ( .I1(n5123), .I2(wb_addr[4]), .O(n4925) );
  ND3S U4146 ( .I1(n4741), .I2(n4740), .I3(n4739), .O(n2593) );
  ND2S U4147 ( .I1(n5123), .I2(wb_addr[3]), .O(n4739) );
  ND2S U4148 ( .I1(n4738), .I2(n5131), .O(n4741) );
  ND3S U4149 ( .I1(n4636), .I2(n4635), .I3(n4634), .O(n2594) );
  ND2S U4150 ( .I1(n5123), .I2(wb_addr[2]), .O(n4634) );
  ND2S U4151 ( .I1(n4596), .I2(n5131), .O(n4636) );
  AO12S U4152 ( .B1(n5113), .B2(n5131), .A1(n5112), .O(n2595) );
  ND3S U4153 ( .I1(n5111), .I2(n5110), .I3(n5109), .O(n5112) );
  AO12S U4154 ( .B1(n5132), .B2(n5131), .A1(n5130), .O(n2596) );
  ND3S U4155 ( .I1(n5129), .I2(n5128), .I3(n5127), .O(n5130) );
  ND2S U4156 ( .I1(n5123), .I2(wb_addr[0]), .O(n5129) );
  ND3S U4157 ( .I1(n3670), .I2(n3669), .I3(n3668), .O(n2597) );
  ND2S U4158 ( .I1(n5092), .I2(n3667), .O(n3668) );
  ND2S U4159 ( .I1(n3655), .I2(n5098), .O(n3670) );
  ND3S U4160 ( .I1(n4367), .I2(n4366), .I3(n4365), .O(n2598) );
  ND3S U4161 ( .I1(n4374), .I2(n4373), .I3(n5109), .O(n2599) );
  AO22S U4162 ( .A1(n3493), .A2(n6298), .B1(n3492), .B2(avg_temp[0]), .O(n2606) );
  AO22S U4163 ( .A1(n3492), .A2(avg_temp[8]), .B1(n3493), .B2(n6269), .O(n2614) );
  ND2S U4164 ( .I1(n5610), .I2(avg_temp[9]), .O(n3671) );
  MUX2S U4165 ( .A(filter_result_reg[24]), .B(filter_result_reg[56]), .S(n6263), .O(n2616) );
  MUX2S U4166 ( .A(filter_result_reg[56]), .B(filter_result_reg[88]), .S(n6263), .O(n2617) );
  MUX2S U4167 ( .A(filter_result_reg[16]), .B(filter_result_reg[48]), .S(n6263), .O(n2618) );
  MUX2S U4168 ( .A(filter_result_reg[48]), .B(filter_result_reg[80]), .S(n6266), .O(n2619) );
  MUX2S U4169 ( .A(filter_result_reg[8]), .B(filter_result_reg[40]), .S(n6266), 
        .O(n2620) );
  MUX2S U4170 ( .A(filter_result_reg[40]), .B(filter_result_reg[72]), .S(n6266), .O(n2621) );
  MUX2S U4171 ( .A(filter_result_reg[0]), .B(filter_result_reg[32]), .S(n6266), 
        .O(n2622) );
  MUX2S U4172 ( .A(filter_result_reg[32]), .B(filter_result_reg[64]), .S(n6266), .O(n2623) );
  MUX2S U4173 ( .A(filter_result_reg[25]), .B(filter_result_reg[57]), .S(n6266), .O(n2625) );
  MUX2S U4174 ( .A(filter_result_reg[57]), .B(filter_result_reg[89]), .S(n6263), .O(n2626) );
  MUX2S U4175 ( .A(filter_result_reg[17]), .B(filter_result_reg[49]), .S(n6263), .O(n2627) );
  MUX2S U4176 ( .A(filter_result_reg[49]), .B(filter_result_reg[81]), .S(n6263), .O(n2628) );
  MUX2S U4177 ( .A(filter_result_reg[9]), .B(filter_result_reg[41]), .S(n6263), 
        .O(n2629) );
  MUX2S U4178 ( .A(filter_result_reg[41]), .B(filter_result_reg[73]), .S(n6263), .O(n2630) );
  MUX2S U4179 ( .A(filter_result_reg[1]), .B(filter_result_reg[33]), .S(n6263), 
        .O(n2631) );
  MUX2S U4180 ( .A(filter_result_reg[33]), .B(filter_result_reg[65]), .S(n6263), .O(n2632) );
  MUX2S U4181 ( .A(filter_result_reg[26]), .B(filter_result_reg[58]), .S(n6263), .O(n2634) );
  MUX2S U4182 ( .A(filter_result_reg[58]), .B(filter_result_reg[90]), .S(n6263), .O(n2635) );
  MUX2S U4183 ( .A(filter_result_reg[18]), .B(filter_result_reg[50]), .S(n6263), .O(n2636) );
  MUX2S U4184 ( .A(filter_result_reg[50]), .B(filter_result_reg[82]), .S(n6263), .O(n2637) );
  MUX2S U4185 ( .A(filter_result_reg[10]), .B(filter_result_reg[42]), .S(n6263), .O(n2638) );
  MUX2S U4186 ( .A(filter_result_reg[42]), .B(filter_result_reg[74]), .S(n6266), .O(n2639) );
  MUX2S U4187 ( .A(filter_result_reg[2]), .B(filter_result_reg[34]), .S(n6266), 
        .O(n2640) );
  MUX2S U4188 ( .A(filter_result_reg[34]), .B(filter_result_reg[66]), .S(n6266), .O(n2641) );
  MUX2S U4189 ( .A(filter_result_reg[27]), .B(filter_result_reg[59]), .S(n6266), .O(n2643) );
  MUX2S U4190 ( .A(filter_result_reg[59]), .B(filter_result_reg[91]), .S(n6263), .O(n2644) );
  MUX2S U4191 ( .A(filter_result_reg[19]), .B(filter_result_reg[51]), .S(n6263), .O(n2645) );
  MUX2S U4192 ( .A(filter_result_reg[51]), .B(filter_result_reg[83]), .S(n6263), .O(n2646) );
  MUX2S U4193 ( .A(filter_result_reg[11]), .B(filter_result_reg[43]), .S(n6263), .O(n2647) );
  MUX2S U4194 ( .A(filter_result_reg[43]), .B(filter_result_reg[75]), .S(n6263), .O(n2648) );
  MUX2S U4195 ( .A(filter_result_reg[3]), .B(filter_result_reg[35]), .S(n6263), 
        .O(n2649) );
  MUX2S U4196 ( .A(filter_result_reg[35]), .B(filter_result_reg[67]), .S(n6266), .O(n2650) );
  MUX2S U4197 ( .A(filter_result_reg[28]), .B(filter_result_reg[60]), .S(n6266), .O(n2652) );
  MUX2S U4198 ( .A(filter_result_reg[60]), .B(filter_result_reg[92]), .S(n6263), .O(n2653) );
  MUX2S U4199 ( .A(filter_result_reg[20]), .B(filter_result_reg[52]), .S(n6266), .O(n2654) );
  MUX2S U4200 ( .A(filter_result_reg[52]), .B(filter_result_reg[84]), .S(n6266), .O(n2655) );
  MUX2S U4201 ( .A(filter_result_reg[12]), .B(filter_result_reg[44]), .S(n6266), .O(n2656) );
  MUX2S U4202 ( .A(filter_result_reg[44]), .B(filter_result_reg[76]), .S(n6266), .O(n2657) );
  MUX2S U4203 ( .A(filter_result_reg[4]), .B(filter_result_reg[36]), .S(n6266), 
        .O(n2658) );
  MUX2S U4204 ( .A(filter_result_reg[36]), .B(filter_result_reg[68]), .S(n6266), .O(n2659) );
  MUX2S U4205 ( .A(filter_result_reg[29]), .B(filter_result_reg[61]), .S(n6266), .O(n2661) );
  MUX2S U4206 ( .A(filter_result_reg[61]), .B(filter_result_reg[93]), .S(n6266), .O(n2662) );
  MUX2S U4207 ( .A(filter_result_reg[21]), .B(filter_result_reg[53]), .S(n6263), .O(n2663) );
  MUX2S U4208 ( .A(filter_result_reg[53]), .B(filter_result_reg[85]), .S(n6263), .O(n2664) );
  MUX2S U4209 ( .A(filter_result_reg[13]), .B(filter_result_reg[45]), .S(n6263), .O(n2665) );
  MUX2S U4210 ( .A(filter_result_reg[45]), .B(filter_result_reg[77]), .S(n6263), .O(n2666) );
  MUX2S U4211 ( .A(filter_result_reg[5]), .B(filter_result_reg[37]), .S(n6263), 
        .O(n2667) );
  MUX2S U4212 ( .A(filter_result_reg[37]), .B(filter_result_reg[69]), .S(n6263), .O(n2668) );
  MUX2S U4213 ( .A(filter_result_reg[30]), .B(filter_result_reg[62]), .S(n6263), .O(n2670) );
  MUX2S U4214 ( .A(filter_result_reg[62]), .B(filter_result_reg[94]), .S(n6263), .O(n2671) );
  MUX2S U4215 ( .A(filter_result_reg[22]), .B(filter_result_reg[54]), .S(n6263), .O(n2672) );
  MUX2S U4216 ( .A(filter_result_reg[54]), .B(filter_result_reg[86]), .S(n6263), .O(n2673) );
  MUX2S U4217 ( .A(filter_result_reg[14]), .B(filter_result_reg[46]), .S(n6263), .O(n2674) );
  MUX2S U4218 ( .A(filter_result_reg[46]), .B(filter_result_reg[78]), .S(n6263), .O(n2675) );
  MUX2S U4219 ( .A(filter_result_reg[6]), .B(filter_result_reg[38]), .S(n6263), 
        .O(n2676) );
  MUX2S U4220 ( .A(filter_result_reg[38]), .B(filter_result_reg[70]), .S(n6263), .O(n2677) );
  MUX2S U4221 ( .A(filter_result_reg[31]), .B(filter_result_reg[63]), .S(n6263), .O(n2704) );
  MUX2S U4222 ( .A(filter_result_reg[63]), .B(filter_result_reg[95]), .S(n6263), .O(n2705) );
  MUX2S U4223 ( .A(filter_result_reg[23]), .B(filter_result_reg[55]), .S(n6263), .O(n2706) );
  MUX2S U4224 ( .A(filter_result_reg[55]), .B(filter_result_reg[87]), .S(n6263), .O(n2707) );
  MUX2S U4225 ( .A(filter_result_reg[15]), .B(filter_result_reg[47]), .S(n6263), .O(n2708) );
  MUX2S U4226 ( .A(filter_result_reg[47]), .B(filter_result_reg[79]), .S(n6263), .O(n2709) );
  MUX2S U4227 ( .A(filter_result_reg[7]), .B(filter_result_reg[39]), .S(n6263), 
        .O(n2710) );
  MUX2S U4228 ( .A(filter_result_reg[39]), .B(filter_result_reg[71]), .S(n6263), .O(n2711) );
  AO22S U4229 ( .A1(n6210), .A2(gray_avg_reg[24]), .B1(n6219), .B2(
        gray_avg_reg[16]), .O(n2760) );
  AO22S U4230 ( .A1(n6210), .A2(gray_avg_reg[25]), .B1(n6219), .B2(
        gray_avg_reg[17]), .O(n2761) );
  AO22S U4231 ( .A1(n6210), .A2(gray_avg_reg[26]), .B1(n6219), .B2(
        gray_avg_reg[18]), .O(n2762) );
  AO22S U4232 ( .A1(n6210), .A2(gray_avg_reg[27]), .B1(n6219), .B2(
        gray_avg_reg[19]), .O(n2763) );
  AO22S U4233 ( .A1(n6210), .A2(gray_avg_reg[28]), .B1(n6219), .B2(
        gray_avg_reg[20]), .O(n2764) );
  AO22S U4234 ( .A1(n6210), .A2(gray_avg_reg[30]), .B1(n6219), .B2(
        gray_avg_reg[22]), .O(n2766) );
  AO22S U4235 ( .A1(n6210), .A2(gray_avg_reg[31]), .B1(n6219), .B2(
        gray_avg_reg[23]), .O(n2767) );
  ND2S U4236 ( .I1(n4876), .I2(n4875), .O(n2768) );
  OR2S U4237 ( .I1(n6219), .I2(n4874), .O(n4875) );
  ND2S U4238 ( .I1(gray_avg_reg[24]), .I2(n6219), .O(n4876) );
  OA12S U4239 ( .B1(n6210), .B2(gray_avg_reg[25]), .A1(n6208), .O(n2769) );
  AO112S U4240 ( .C1(avg_temp[1]), .C2(n6207), .A1(n6206), .B1(n6219), .O(
        n6208) );
  OA12S U4241 ( .B1(n6204), .B2(n6293), .A1(n6203), .O(n6205) );
  ND2S U4242 ( .I1(n6210), .I2(n6199), .O(n6200) );
  AO22S U4243 ( .A1(n6196), .A2(gray_max_temp[31]), .B1(n6193), .B2(
        gray_max_temp[23]), .O(n2778) );
  AO22S U4244 ( .A1(n6196), .A2(gray_max_temp[29]), .B1(n6188), .B2(
        gray_max_temp[21]), .O(n2782) );
  AO22S U4245 ( .A1(n6196), .A2(gray_max_temp[28]), .B1(n6177), .B2(
        gray_max_temp[20]), .O(n2786) );
  AO22S U4246 ( .A1(n6196), .A2(gray_max_temp[27]), .B1(n6193), .B2(
        gray_max_temp[19]), .O(n2790) );
  AO22S U4247 ( .A1(n6196), .A2(gray_max_temp[26]), .B1(n6193), .B2(
        gray_max_temp[18]), .O(n2794) );
  AO22S U4248 ( .A1(n6196), .A2(gray_max_temp[25]), .B1(n6188), .B2(
        gray_max_temp[17]), .O(n2798) );
  AO22S U4249 ( .A1(n6196), .A2(gray_max_temp[24]), .B1(n6177), .B2(
        gray_max_temp[16]), .O(n2802) );
  AO22S U4250 ( .A1(n6196), .A2(gray_max_temp[30]), .B1(n6188), .B2(
        gray_max_temp[22]), .O(n2806) );
  AO222S U4251 ( .A1(n5473), .A2(find_median_inst_mid_mid_reg[0]), .B1(n5472), 
        .B2(find_median_inst_max_min_reg[0]), .C1(n5474), .C2(
        find_median_inst_min_pool_temp[0]), .O(find_median_inst_final_mid[0])
         );
  AO222S U4252 ( .A1(n5389), .A2(find_median_inst_mid2_reg[0]), .B1(n5388), 
        .B2(find_median_inst_mid1_reg[0]), .C1(n5390), .C2(
        find_median_inst_mid3_reg[0]), .O(find_median_inst_mid_mid[0]) );
  AO222S U4253 ( .A1(n5474), .A2(find_median_inst_min_pool_temp[1]), .B1(
        find_median_inst_mid_mid_reg[1]), .B2(n5473), .C1(
        find_median_inst_max_min_reg[1]), .C2(n5472), .O(
        find_median_inst_final_mid[1]) );
  AO222S U4254 ( .A1(n5389), .A2(find_median_inst_mid2_reg[1]), .B1(n5388), 
        .B2(find_median_inst_mid1_reg[1]), .C1(n5390), .C2(
        find_median_inst_mid3_reg[1]), .O(find_median_inst_mid_mid[1]) );
  AO222S U4255 ( .A1(n5474), .A2(find_median_inst_min_pool_temp[4]), .B1(
        find_median_inst_mid_mid_reg[4]), .B2(n5473), .C1(
        find_median_inst_max_min_reg[4]), .C2(n5472), .O(
        find_median_inst_final_mid[4]) );
  AO222S U4256 ( .A1(n5390), .A2(find_median_inst_mid3_reg[4]), .B1(
        find_median_inst_mid1_reg[4]), .B2(n5388), .C1(
        find_median_inst_mid2_reg[4]), .C2(n5389), .O(
        find_median_inst_mid_mid[4]) );
  AO222S U4257 ( .A1(n5390), .A2(find_median_inst_mid3_reg[7]), .B1(
        find_median_inst_mid2_reg[7]), .B2(n5389), .C1(
        find_median_inst_mid1_reg[7]), .C2(n5388), .O(
        find_median_inst_mid_mid[7]) );
  AO222S U4258 ( .A1(n5474), .A2(find_median_inst_min_pool_temp[7]), .B1(
        find_median_inst_mid_mid_reg[7]), .B2(n5473), .C1(
        find_median_inst_max_min_reg[7]), .C2(n5472), .O(
        find_median_inst_final_mid[7]) );
  MOAI1S U4259 ( .A1(n4782), .A2(n61290), .B1(n4956), .B2(conv_temp[17]), .O(
        n2866) );
  MOAI1S U4260 ( .A1(n4782), .A2(n61300), .B1(n4956), .B2(conv_temp[16]), .O(
        n2867) );
  MUX2S U4261 ( .A(n5063), .B(n5064), .S(wb_addr[0]), .O(n3204) );
  MUX2S U4262 ( .A(n5014), .B(n5016), .S(wb_addr[7]), .O(n3205) );
  AN2S U4263 ( .I1(n5012), .I2(n5063), .O(n5014) );
  ND3S U4264 ( .I1(n4632), .I2(n3532), .I3(n3531), .O(n6300) );
  ND3S U4265 ( .I1(n3529), .I2(n5984), .I3(n3528), .O(n3532) );
  MUX2S U4266 ( .A(n5715), .B(n5695), .S(cal_count_10[0]), .O(n3217) );
  INV1S U4267 ( .I(n5695), .O(n6301) );
  ND3S U4268 ( .I1(n4985), .I2(n4184), .I3(n4183), .O(n3404) );
  AO22S U4269 ( .A1(n5626), .A2(wgt_temp[6]), .B1(n5625), .B2(n5624), .O(n3347) );
  AO222S U4270 ( .A1(n5626), .A2(wgt_temp[5]), .B1(n5624), .B2(n5622), .C1(
        image[7]), .C2(n5621), .O(n3348) );
  AO222S U4271 ( .A1(n5626), .A2(wgt_temp[4]), .B1(n5624), .B2(n5619), .C1(
        image[6]), .C2(n5621), .O(n3349) );
  AO222S U4272 ( .A1(n5626), .A2(wgt_temp[3]), .B1(n5624), .B2(n5617), .C1(
        image[5]), .C2(n5621), .O(n3350) );
  AO222S U4273 ( .A1(n5626), .A2(wgt_temp[2]), .B1(n5624), .B2(n5615), .C1(
        image[4]), .C2(n5621), .O(n3351) );
  AO222S U4274 ( .A1(n5626), .A2(wgt_temp[1]), .B1(n5624), .B2(n5613), .C1(
        image[3]), .C2(n5621), .O(n3352) );
  AO222S U4275 ( .A1(n5626), .A2(wgt_temp[0]), .B1(n5611), .B2(n5624), .C1(
        image[2]), .C2(n5621), .O(n3353) );
  XNR2HS U4276 ( .I1(wgt_temp[7]), .I2(n3674), .O(n3678) );
  MOAI1S U4277 ( .A1(n5608), .A2(n3900), .B1(max_temp[6]), .B2(n5607), .O(
        n3362) );
  AO12S U4278 ( .B1(action_idx[3]), .B2(n5569), .A1(n5570), .O(n3395) );
  OA12S U4279 ( .B1(action_idx[2]), .B2(n5579), .A1(n5569), .O(n3396) );
  AO222S U4280 ( .A1(n3647), .A2(filter_result_reg[8]), .B1(pool_temp[8]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[8]), .O(n2900) );
  AO222S U4281 ( .A1(n3647), .A2(filter_result_reg[24]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[24]), .C1(pool_temp[24]), .C2(n6056), .O(n2916)
         );
  AO222S U4282 ( .A1(n3647), .A2(filter_result_reg[16]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[16]), .C1(pool_temp[16]), .C2(n6056), .O(n3089)
         );
  AO222S U4283 ( .A1(n3647), .A2(filter_result_reg[0]), .B1(pool_temp[0]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[0]), .O(n3073) );
  ND3S U4284 ( .I1(n4503), .I2(n4502), .I3(n4501), .O(n3001) );
  AO222S U4285 ( .A1(n5932), .A2(SRAM_out_buffer[24]), .B1(n5964), .B2(n5931), 
        .C1(n5930), .C2(SRAM_out_buffer[56]), .O(n3002) );
  AO222S U4286 ( .A1(n6064), .A2(median_in[56]), .B1(n5939), .B2(median_in[48]), .C1(n4935), .C2(SRAM_out_buffer[88]), .O(n3004) );
  ND2S U4287 ( .I1(n4916), .I2(n4915), .O(n3006) );
  OR3S U4288 ( .I1(n4919), .I2(n4918), .I3(n4917), .O(n6305) );
  ND3S U4289 ( .I1(n4704), .I2(n4703), .I3(n4702), .O(n3008) );
  ND3S U4290 ( .I1(n4719), .I2(n4718), .I3(n4717), .O(n3053) );
  ND2S U4291 ( .I1(SRAM_out_buffer[48]), .I2(n4772), .O(n4717) );
  ND3S U4292 ( .I1(n4469), .I2(n4468), .I3(n4467), .O(n3133) );
  AO222S U4293 ( .A1(n5765), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[0]), 
        .C1(n5930), .C2(SRAM_out_buffer[32]), .O(n3160) );
  ND2S U4294 ( .I1(n4907), .I2(n4906), .O(n3055) );
  AO222S U4295 ( .A1(n5773), .A2(SRAM_out_buffer[64]), .B1(n4385), .B2(
        window_0__4__0_), .C1(n5771), .C2(SRAM_out_buffer[72]), .O(n3135) );
  ND3S U4296 ( .I1(n4707), .I2(n4706), .I3(n4705), .O(n3056) );
  ND3S U4297 ( .I1(n4400), .I2(n4399), .I3(n4398), .O(n3136) );
  AO222S U4298 ( .A1(n3647), .A2(filter_result_reg[9]), .B1(pool_temp[9]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[9]), .O(n2898) );
  AO222S U4299 ( .A1(n3647), .A2(filter_result_reg[25]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[25]), .C1(pool_temp[25]), .C2(n6056), .O(n2914)
         );
  AO222S U4300 ( .A1(n3647), .A2(filter_result_reg[17]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[17]), .C1(pool_temp[17]), .C2(n6056), .O(n3087)
         );
  AO222S U4301 ( .A1(n3647), .A2(filter_result_reg[1]), .B1(pool_temp[1]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[1]), .O(n3071) );
  AO12S U4302 ( .B1(n4978), .B2(n3517), .A1(n4977), .O(n2987) );
  ND3S U4303 ( .I1(n4976), .I2(n4975), .I3(n4974), .O(n4977) );
  ND2S U4304 ( .I1(n4981), .I2(median_in[9]), .O(n4976) );
  OR3B2S U4305 ( .I1(n4978), .B1(n4449), .B2(n4975), .O(n2988) );
  AO222S U4306 ( .A1(n6064), .A2(median_in[57]), .B1(n5939), .B2(median_in[49]), .C1(SRAM_out_buffer[89]), .C2(n4935), .O(n2992) );
  ND2S U4307 ( .I1(n4901), .I2(n4900), .O(n2993) );
  ND2S U4308 ( .I1(n4865), .I2(n4864), .O(n2994) );
  AO112S U4309 ( .C1(median_in[25]), .C2(n5939), .A1(n4941), .B1(n4940), .O(
        n2995) );
  ND3S U4310 ( .I1(n4759), .I2(n4758), .I3(n4757), .O(n3047) );
  ND3S U4311 ( .I1(n4507), .I2(n4506), .I3(n4505), .O(n3127) );
  AO222S U4312 ( .A1(n5807), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[1]), 
        .C1(n5930), .C2(SRAM_out_buffer[33]), .O(n3157) );
  ND2S U4313 ( .I1(n4888), .I2(n4887), .O(n3049) );
  AO222S U4314 ( .A1(n4385), .A2(window_0__4__1_), .B1(n5773), .B2(
        SRAM_out_buffer[65]), .C1(n5771), .C2(SRAM_out_buffer[73]), .O(n3129)
         );
  ND3S U4315 ( .I1(n4669), .I2(n4668), .I3(n4667), .O(n3050) );
  ND3S U4316 ( .I1(n4397), .I2(n4396), .I3(n4395), .O(n3130) );
  AO222S U4317 ( .A1(n3647), .A2(filter_result_reg[10]), .B1(pool_temp[10]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[10]), .O(n2896) );
  AO222S U4318 ( .A1(n3647), .A2(filter_result_reg[26]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[26]), .C1(pool_temp[26]), .C2(n6056), .O(n2912)
         );
  AO222S U4319 ( .A1(n3647), .A2(filter_result_reg[18]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[18]), .C1(pool_temp[18]), .C2(n6056), .O(n3085)
         );
  AO222S U4320 ( .A1(n3647), .A2(filter_result_reg[2]), .B1(pool_temp[2]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[2]), .O(n3069) );
  ND3S U4321 ( .I1(n4444), .I2(n4443), .I3(n4442), .O(n2975) );
  OA22S U4322 ( .A1(n5265), .A2(n6068), .B1(n5918), .B2(n4441), .O(n4443) );
  ND3S U4323 ( .I1(n4441), .I2(n4431), .I3(n4442), .O(n2976) );
  ND3S U4324 ( .I1(n4724), .I2(n4723), .I3(n4722), .O(n3041) );
  ND2S U4325 ( .I1(n4767), .I2(SRAM_out_buffer[42]), .O(n4722) );
  AO222S U4326 ( .A1(n5886), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[18]), 
        .C1(SRAM_out_buffer[50]), .C2(n5930), .O(n3042) );
  ND3S U4327 ( .I1(n4518), .I2(n4517), .I3(n4516), .O(n2981) );
  ND2S U4328 ( .I1(n4889), .I2(window_0__3__2_), .O(n4517) );
  AO112S U4329 ( .C1(median_in[26]), .C2(n5939), .A1(n4970), .B1(n4939), .O(
        n2983) );
  ND2S U4330 ( .I1(n4891), .I2(n4890), .O(n3043) );
  ND3S U4331 ( .I1(n4678), .I2(n4677), .I3(n4676), .O(n3044) );
  AO222S U4332 ( .A1(n5800), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[10]), 
        .C1(SRAM_out_buffer[42]), .C2(n5916), .O(n3122) );
  AO222S U4333 ( .A1(n4385), .A2(window_0__4__2_), .B1(n5773), .B2(
        SRAM_out_buffer[66]), .C1(n5771), .C2(SRAM_out_buffer[74]), .O(n3123)
         );
  ND3S U4334 ( .I1(n4403), .I2(n4402), .I3(n4401), .O(n3124) );
  AO222S U4335 ( .A1(n3647), .A2(filter_result_reg[11]), .B1(pool_temp[11]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[11]), .O(n2894) );
  AO222S U4336 ( .A1(n3647), .A2(filter_result_reg[27]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[27]), .C1(pool_temp[27]), .C2(n6056), .O(n2910)
         );
  AO222S U4337 ( .A1(n3647), .A2(filter_result_reg[19]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[19]), .C1(pool_temp[19]), .C2(n6056), .O(n3083)
         );
  AO222S U4338 ( .A1(n3647), .A2(filter_result_reg[3]), .B1(pool_temp[3]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[3]), .O(n3067) );
  ND2S U4339 ( .I1(n4980), .I2(n4895), .O(n2964) );
  ND3S U4340 ( .I1(n4779), .I2(n4778), .I3(n4777), .O(n3035) );
  ND2S U4341 ( .I1(n4889), .I2(window_2__4__3_), .O(n4777) );
  AO222S U4342 ( .A1(n5887), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[19]), 
        .C1(SRAM_out_buffer[51]), .C2(n5916), .O(n3036) );
  ND2S U4343 ( .I1(n4897), .I2(n4896), .O(n2969) );
  ND2S U4344 ( .I1(n4860), .I2(n4859), .O(n2970) );
  AO112S U4345 ( .C1(median_in[27]), .C2(n5939), .A1(n5892), .B1(n5891), .O(
        n2971) );
  ND2S U4346 ( .I1(n4886), .I2(n4885), .O(n3037) );
  ND3S U4347 ( .I1(n4666), .I2(n4665), .I3(n4664), .O(n3038) );
  AO222S U4348 ( .A1(n5797), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[11]), 
        .C1(SRAM_out_buffer[43]), .C2(n5916), .O(n3116) );
  AO222S U4349 ( .A1(n4385), .A2(window_0__4__3_), .B1(n5773), .B2(
        SRAM_out_buffer[67]), .C1(n5771), .C2(SRAM_out_buffer[75]), .O(n3117)
         );
  ND3S U4350 ( .I1(n4412), .I2(n4411), .I3(n4410), .O(n3118) );
  AO222S U4351 ( .A1(n3647), .A2(filter_result_reg[12]), .B1(pool_temp[12]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[12]), .O(n2892) );
  AO222S U4352 ( .A1(n3647), .A2(filter_result_reg[28]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[28]), .C1(pool_temp[28]), .C2(n6056), .O(n2908)
         );
  AO222S U4353 ( .A1(n3647), .A2(filter_result_reg[20]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[20]), .C1(pool_temp[20]), .C2(n6056), .O(n3081)
         );
  AO222S U4354 ( .A1(n3647), .A2(filter_result_reg[4]), .B1(pool_temp[4]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[4]), .O(n3065) );
  OA22S U4355 ( .A1(n5906), .A2(n6068), .B1(n5918), .B2(n5905), .O(n5908) );
  ND3S U4356 ( .I1(n5905), .I2(n4110), .I3(n5907), .O(n2952) );
  ND3S U4357 ( .I1(n4770), .I2(n4769), .I3(n4768), .O(n3029) );
  AO222S U4358 ( .A1(n5951), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[20]), 
        .C1(SRAM_out_buffer[52]), .C2(n5916), .O(n3030) );
  ND2S U4359 ( .I1(n4899), .I2(n4898), .O(n2957) );
  ND2S U4360 ( .I1(n4863), .I2(n4862), .O(n2958) );
  AO112S U4361 ( .C1(median_in[28]), .C2(n5939), .A1(n5901), .B1(n5900), .O(
        n2959) );
  ND2S U4362 ( .I1(n4909), .I2(n4908), .O(n3031) );
  ND3S U4363 ( .I1(n4672), .I2(n4671), .I3(n4670), .O(n3032) );
  AO222S U4364 ( .A1(n5798), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[12]), 
        .C1(SRAM_out_buffer[44]), .C2(n5916), .O(n3110) );
  AO222S U4365 ( .A1(n4385), .A2(window_0__4__4_), .B1(n5773), .B2(
        SRAM_out_buffer[68]), .C1(n5771), .C2(SRAM_out_buffer[76]), .O(n3111)
         );
  ND3S U4366 ( .I1(n4409), .I2(n4408), .I3(n4407), .O(n3112) );
  AO222S U4367 ( .A1(n3647), .A2(filter_result_reg[13]), .B1(pool_temp[13]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[13]), .O(n2890) );
  AO222S U4368 ( .A1(n3647), .A2(filter_result_reg[29]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[29]), .C1(pool_temp[29]), .C2(n6056), .O(n2906)
         );
  AO222S U4369 ( .A1(n3647), .A2(filter_result_reg[21]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[21]), .C1(pool_temp[21]), .C2(n6056), .O(n3079)
         );
  AO222S U4370 ( .A1(n3647), .A2(filter_result_reg[5]), .B1(pool_temp[5]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[5]), .O(n3063) );
  OA22S U4371 ( .A1(n5919), .A2(n5942), .B1(n5918), .B2(n5917), .O(n5921) );
  ND3S U4372 ( .I1(n5917), .I2(n4423), .I3(n5920), .O(n2940) );
  ND3S U4373 ( .I1(n4754), .I2(n4753), .I3(n4752), .O(n2941) );
  OA12S U4374 ( .B1(n5942), .B2(n5269), .A1(n4750), .O(n4753) );
  ND3S U4375 ( .I1(n4764), .I2(n4763), .I3(n4762), .O(n3023) );
  AO222S U4376 ( .A1(n5948), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[21]), 
        .C1(SRAM_out_buffer[53]), .C2(n5916), .O(n3024) );
  ND2S U4377 ( .I1(n4913), .I2(n4912), .O(n2946) );
  AO112S U4378 ( .C1(median_in[29]), .C2(n5939), .A1(n5912), .B1(n5911), .O(
        n2947) );
  ND3S U4379 ( .I1(n4712), .I2(n4711), .I3(n4710), .O(n2948) );
  ND2S U4380 ( .I1(n4905), .I2(n4904), .O(n3025) );
  ND3S U4381 ( .I1(n4496), .I2(n4495), .I3(n4494), .O(n3103) );
  AO222S U4382 ( .A1(n5792), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[13]), 
        .C1(SRAM_out_buffer[45]), .C2(n5930), .O(n3104) );
  AO222S U4383 ( .A1(n4385), .A2(window_0__4__5_), .B1(n5773), .B2(
        SRAM_out_buffer[69]), .C1(n5771), .C2(SRAM_out_buffer[77]), .O(n3105)
         );
  ND3S U4384 ( .I1(n4406), .I2(n4405), .I3(n4404), .O(n3106) );
  AO222S U4385 ( .A1(n3647), .A2(filter_result_reg[14]), .B1(pool_temp[14]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[14]), .O(n2888) );
  AO222S U4386 ( .A1(n3647), .A2(filter_result_reg[30]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[30]), .C1(pool_temp[30]), .C2(n6056), .O(n2904)
         );
  AO222S U4387 ( .A1(n3647), .A2(filter_result_reg[22]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[22]), .C1(pool_temp[22]), .C2(n6056), .O(n3077)
         );
  AO222S U4388 ( .A1(n3647), .A2(filter_result_reg[6]), .B1(pool_temp[6]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[6]), .O(n3061) );
  ND3S U4389 ( .I1(n4440), .I2(n4439), .I3(n4438), .O(n2927) );
  OA22S U4390 ( .A1(n5270), .A2(n6068), .B1(n5918), .B2(n4437), .O(n4439) );
  ND3S U4391 ( .I1(n4437), .I2(n4427), .I3(n4438), .O(n2928) );
  ND3S U4392 ( .I1(n4729), .I2(n4728), .I3(n4727), .O(n3017) );
  AO222S U4393 ( .A1(n5949), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[22]), 
        .C1(SRAM_out_buffer[54]), .C2(n5916), .O(n3018) );
  ND2S U4394 ( .I1(n4878), .I2(n4877), .O(n2933) );
  ND2S U4395 ( .I1(n4911), .I2(n4910), .O(n2934) );
  AO112S U4396 ( .C1(median_in[30]), .C2(n5939), .A1(n5925), .B1(n5924), .O(
        n2935) );
  ND2S U4397 ( .I1(n4882), .I2(n4881), .O(n3019) );
  ND3S U4398 ( .I1(n4681), .I2(n4680), .I3(n4679), .O(n3020) );
  ND3S U4399 ( .I1(n4490), .I2(n4489), .I3(n4488), .O(n3097) );
  AO222S U4400 ( .A1(n5772), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[14]), 
        .C1(SRAM_out_buffer[46]), .C2(n5930), .O(n3098) );
  AO222S U4401 ( .A1(n4385), .A2(window_0__4__6_), .B1(n5773), .B2(
        SRAM_out_buffer[70]), .C1(n5771), .C2(SRAM_out_buffer[78]), .O(n3099)
         );
  ND3S U4402 ( .I1(n4415), .I2(n4414), .I3(n4413), .O(n3100) );
  OR3B2S U4403 ( .I1(n6063), .B1(n4453), .B2(n6065), .O(n2885) );
  ND3S U4404 ( .I1(n4686), .I2(n4685), .I3(n4684), .O(n2886) );
  AO222S U4405 ( .A1(n3647), .A2(filter_result_reg[15]), .B1(pool_temp[15]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[15]), .O(n2902) );
  ND3S U4406 ( .I1(n4734), .I2(n4733), .I3(n4732), .O(n3011) );
  ND2S U4407 ( .I1(SRAM_out_buffer[55]), .I2(n4772), .O(n4732) );
  AO222S U4408 ( .A1(n5969), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[23]), 
        .C1(SRAM_out_buffer[55]), .C2(n5916), .O(n3012) );
  ND2S U4409 ( .I1(n4880), .I2(n4879), .O(n2921) );
  ND2S U4410 ( .I1(n4867), .I2(n4866), .O(n2922) );
  AO112S U4411 ( .C1(median_in[31]), .C2(n5939), .A1(n5938), .B1(n5937), .O(
        n2923) );
  ND3S U4412 ( .I1(n4660), .I2(n4659), .I3(n4658), .O(n2924) );
  ND2S U4413 ( .I1(n4884), .I2(n4883), .O(n3013) );
  ND3S U4414 ( .I1(n4663), .I2(n4662), .I3(n4661), .O(n3014) );
  AO222S U4415 ( .A1(n5884), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[15]), 
        .C1(SRAM_out_buffer[47]), .C2(n5930), .O(n3060) );
  AO222S U4416 ( .A1(n3647), .A2(filter_result_reg[7]), .B1(pool_temp[7]), 
        .B2(n6056), .C1(n6055), .C2(SRAM_64X32_in_decode[7]), .O(n3075) );
  AO222S U4417 ( .A1(n3647), .A2(filter_result_reg[23]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[23]), .C1(pool_temp[23]), .C2(n6056), .O(n3091)
         );
  AO222S U4418 ( .A1(n4385), .A2(window_0__4__7_), .B1(n5773), .B2(
        SRAM_out_buffer[71]), .C1(n5771), .C2(SRAM_out_buffer[79]), .O(n3093)
         );
  ND3S U4419 ( .I1(n4419), .I2(n4418), .I3(n4417), .O(n3094) );
  AO222S U4420 ( .A1(n5885), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[16]), 
        .C1(SRAM_out_buffer[48]), .C2(n5916), .O(n3054) );
  AO222S U4421 ( .A1(n5805), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[8]), 
        .C1(SRAM_out_buffer[40]), .C2(n5916), .O(n3134) );
  AO222S U4422 ( .A1(n5960), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[17]), 
        .C1(SRAM_out_buffer[49]), .C2(n5930), .O(n3048) );
  AO222S U4423 ( .A1(n5804), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[9]), 
        .C1(SRAM_out_buffer[41]), .C2(n5916), .O(n3128) );
  AO222S U4424 ( .A1(n5932), .A2(SRAM_out_buffer[26]), .B1(n5961), .B2(n5931), 
        .C1(n5930), .C2(SRAM_out_buffer[58]), .O(n2978) );
  AO222S U4425 ( .A1(n5806), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[2]), 
        .C1(n5930), .C2(SRAM_out_buffer[34]), .O(n3154) );
  AO222S U4426 ( .A1(n5799), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[3]), 
        .C1(n5930), .C2(SRAM_out_buffer[35]), .O(n3151) );
  AO222S U4427 ( .A1(n5932), .A2(SRAM_out_buffer[28]), .B1(n5955), .B2(n5931), 
        .C1(n5930), .C2(SRAM_out_buffer[60]), .O(n2954) );
  AO222S U4428 ( .A1(n5793), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[4]), 
        .C1(n5930), .C2(SRAM_out_buffer[36]), .O(n3148) );
  AO222S U4429 ( .A1(n5932), .A2(SRAM_out_buffer[29]), .B1(n5950), .B2(n5931), 
        .C1(n5916), .C2(SRAM_out_buffer[61]), .O(n2942) );
  AO222S U4430 ( .A1(n5791), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[5]), 
        .C1(n5930), .C2(SRAM_out_buffer[37]), .O(n3145) );
  AO222S U4431 ( .A1(n5932), .A2(SRAM_out_buffer[30]), .B1(n5967), .B2(n5931), 
        .C1(n5930), .C2(SRAM_out_buffer[62]), .O(n2930) );
  AO222S U4432 ( .A1(n5813), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[6]), 
        .C1(n5930), .C2(SRAM_out_buffer[38]), .O(n3142) );
  AO222S U4433 ( .A1(n5850), .A2(n5931), .B1(n5932), .B2(SRAM_out_buffer[7]), 
        .C1(n5930), .C2(SRAM_out_buffer[39]), .O(n3139) );
  AO222S U4434 ( .A1(n3647), .A2(filter_result_reg[31]), .B1(n6055), .B2(
        SRAM_64X32_in_decode[31]), .C1(pool_temp[31]), .C2(n6056), .O(n3163)
         );
  MUX2S U4435 ( .A(action[1]), .B(action_reg_0__1_), .S(n4989), .O(n3372) );
  MUX2S U4436 ( .A(action[0]), .B(action_reg_0__0_), .S(n4989), .O(n3373) );
  HA1S U4437 ( .A(n3972), .B(n3971), .C(n3969), .S(N6116) );
  XOR3S U4438 ( .I1(n3980), .I2(n3979), .I3(mult_x_231_n11), .O(N6123) );
  MUX2S U4439 ( .A(template[1]), .B(template_reg[65]), .S(n61240), .O(n3271)
         );
  MUX2S U4440 ( .A(template[2]), .B(template_reg[66]), .S(n61240), .O(n3272)
         );
  MUX2S U4441 ( .A(template[3]), .B(template_reg[67]), .S(n61240), .O(n3273)
         );
  MUX2S U4442 ( .A(template[4]), .B(template_reg[68]), .S(n61240), .O(n3274)
         );
  MUX2S U4443 ( .A(template[0]), .B(template_reg[64]), .S(n61240), .O(n3278)
         );
  MUX2S U4444 ( .A(template[1]), .B(template_reg[1]), .S(n5637), .O(n3335) );
  MUX2S U4445 ( .A(template[2]), .B(template_reg[2]), .S(n5637), .O(n3336) );
  MUX2S U4446 ( .A(template[3]), .B(template_reg[3]), .S(n5637), .O(n3337) );
  MUX2S U4447 ( .A(template[4]), .B(template_reg[4]), .S(n5637), .O(n3338) );
  MUX2S U4448 ( .A(template[0]), .B(template_reg[0]), .S(n5637), .O(n3342) );
  MUX2S U4449 ( .A(template[1]), .B(template_reg[49]), .S(n5643), .O(n3287) );
  MUX2S U4450 ( .A(template[2]), .B(template_reg[50]), .S(n5643), .O(n3288) );
  MUX2S U4451 ( .A(template[3]), .B(template_reg[51]), .S(n5643), .O(n3289) );
  MUX2S U4452 ( .A(template[4]), .B(template_reg[52]), .S(n5643), .O(n3290) );
  MUX2S U4453 ( .A(template[0]), .B(template_reg[48]), .S(n5643), .O(n3294) );
  MUX2S U4454 ( .A(template[1]), .B(template_reg[33]), .S(n5641), .O(n3303) );
  MUX2S U4455 ( .A(template[2]), .B(template_reg[34]), .S(n5641), .O(n3304) );
  MUX2S U4456 ( .A(template[3]), .B(template_reg[35]), .S(n5641), .O(n3305) );
  MUX2S U4457 ( .A(template[4]), .B(template_reg[36]), .S(n5641), .O(n3306) );
  MUX2S U4458 ( .A(template[0]), .B(template_reg[32]), .S(n5641), .O(n3310) );
  MUX2S U4459 ( .A(template[1]), .B(template_reg[17]), .S(n5639), .O(n3319) );
  MUX2S U4460 ( .A(template[2]), .B(template_reg[18]), .S(n5639), .O(n3320) );
  MUX2S U4461 ( .A(template[3]), .B(template_reg[19]), .S(n5639), .O(n3321) );
  MUX2S U4462 ( .A(template[4]), .B(template_reg[20]), .S(n5639), .O(n3322) );
  MUX2S U4463 ( .A(template[0]), .B(template_reg[16]), .S(n5639), .O(n3326) );
  MUX2S U4464 ( .A(template[1]), .B(template_reg[57]), .S(n5644), .O(n3279) );
  MUX2S U4465 ( .A(template[2]), .B(template_reg[58]), .S(n5644), .O(n3280) );
  MUX2S U4466 ( .A(template[3]), .B(template_reg[59]), .S(n5644), .O(n3281) );
  MUX2S U4467 ( .A(template[4]), .B(template_reg[60]), .S(n5644), .O(n3282) );
  MUX2S U4468 ( .A(template[0]), .B(template_reg[56]), .S(n5644), .O(n3286) );
  MUX2S U4469 ( .A(template[1]), .B(template_reg[25]), .S(n5640), .O(n3311) );
  MUX2S U4470 ( .A(template[2]), .B(template_reg[26]), .S(n5640), .O(n3312) );
  MUX2S U4471 ( .A(template[3]), .B(template_reg[27]), .S(n5640), .O(n3313) );
  MUX2S U4472 ( .A(template[4]), .B(template_reg[28]), .S(n5640), .O(n3314) );
  MUX2S U4473 ( .A(template[0]), .B(template_reg[24]), .S(n5640), .O(n3318) );
  MUX2S U4474 ( .A(template[1]), .B(template_reg[41]), .S(n5642), .O(n3295) );
  MUX2S U4475 ( .A(template[2]), .B(template_reg[42]), .S(n5642), .O(n3296) );
  MUX2S U4476 ( .A(template[3]), .B(template_reg[43]), .S(n5642), .O(n3297) );
  MUX2S U4477 ( .A(template[4]), .B(template_reg[44]), .S(n5642), .O(n3298) );
  MUX2S U4478 ( .A(template[0]), .B(template_reg[40]), .S(n5642), .O(n3302) );
  MUX2S U4479 ( .A(template[1]), .B(template_reg[9]), .S(n5638), .O(n3327) );
  MUX2S U4480 ( .A(template[2]), .B(template_reg[10]), .S(n5638), .O(n3328) );
  MUX2S U4481 ( .A(template[3]), .B(template_reg[11]), .S(n5638), .O(n3329) );
  MUX2S U4482 ( .A(template[4]), .B(template_reg[12]), .S(n5638), .O(n3330) );
  MUX2S U4483 ( .A(template[0]), .B(template_reg[8]), .S(n5638), .O(n3334) );
  NR2T U4484 ( .I1(n4082), .I2(n5668), .O(n4193) );
  MXL2HS U4485 ( .A(mult_x_231_n8), .B(mult_x_231_n7), .S(mult_x_231_n11), 
        .OB(n3901) );
  ND3 U4486 ( .I1(n4920), .I2(n6069), .I3(n5918), .O(n3491) );
  INV1S U4487 ( .I(n3492), .O(n3493) );
  BUF2 U4488 ( .I(rst_n), .O(n6308) );
  AOI112HS U4489 ( .C1(template_reg[8]), .C2(n3806), .A1(n3746), .B1(n3745), 
        .O(n3494) );
  AOI112HS U4490 ( .C1(n3806), .C2(template_reg[15]), .A1(n3792), .B1(n3791), 
        .O(n3495) );
  AOI112HS U4491 ( .C1(template_reg[11]), .C2(n3806), .A1(n3711), .B1(n3710), 
        .O(n3496) );
  AOI112HS U4492 ( .C1(template_reg[10]), .C2(n3806), .A1(n3757), .B1(n3756), 
        .O(n3499) );
  AOI112HS U4493 ( .C1(n3806), .C2(template_reg[14]), .A1(n3766), .B1(n3765), 
        .O(n3500) );
  NR2P U4494 ( .I1(n4599), .I2(n5759), .O(n5942) );
  AOI112HS U4495 ( .C1(template_reg[9]), .C2(n3806), .A1(n3735), .B1(n3734), 
        .O(n3501) );
  AOI112HS U4496 ( .C1(n3806), .C2(template_reg[13]), .A1(n3698), .B1(n3697), 
        .O(n3502) );
  AOI112HS U4497 ( .C1(template_reg[12]), .C2(n3806), .A1(n3722), .B1(n3721), 
        .O(n3503) );
  XOR2HS U4498 ( .I1(n4120), .I2(n4119), .O(n3504) );
  INV2 U4499 ( .I(n4432), .O(n4889) );
  NR2 U4500 ( .I1(n5751), .I2(n5077), .O(n3506) );
  OA12S U4501 ( .B1(n3577), .B2(n3576), .A1(n3575), .O(n3507) );
  INV1S U4502 ( .I(n4569), .O(n3550) );
  NR2T U4503 ( .I1(n4067), .I2(n3993), .O(n3537) );
  INV1S U4504 ( .I(n3517), .O(n5918) );
  AOI112HS U4505 ( .C1(n3806), .C2(median_in[15]), .A1(n3805), .B1(n3804), .O(
        n3509) );
  AOI112HS U4506 ( .C1(n3806), .C2(median_in[13]), .A1(n3740), .B1(n3739), .O(
        n3510) );
  AN3 U4507 ( .I1(n3705), .I2(n3704), .I3(n3703), .O(n3511) );
  AOI112HS U4508 ( .C1(n3806), .C2(median_in[10]), .A1(n3716), .B1(n3715), .O(
        n3512) );
  MAO222 U4509 ( .A1(pool_temp[31]), .B1(n6029), .C1(n5991), .O(n5992) );
  MAO222 U4510 ( .A1(pool_temp[6]), .B1(n5881), .C1(n5847), .O(n5848) );
  AOI112HS U4511 ( .C1(median_in[8]), .C2(n3806), .A1(n3751), .B1(n3750), .O(
        n3515) );
  NR2 U4512 ( .I1(max_temp[2]), .I2(n5603), .O(n3891) );
  ND3S U4513 ( .I1(n6089), .I2(n6088), .I3(wait_conv_out_count[0]), .O(n6099)
         );
  ND3S U4514 ( .I1(n3648), .I2(n3647), .I3(n4988), .O(n3656) );
  MAO222 U4515 ( .A1(pool_temp[13]), .B1(n6046), .C1(n6021), .O(n6022) );
  ND3S U4516 ( .I1(n5803), .I2(n5802), .I3(n5801), .O(n5833) );
  ND3S U4517 ( .I1(n6110), .I2(n6109), .I3(n6108), .O(n6111) );
  ND2 U4518 ( .I1(n4620), .I2(n4539), .O(n4562) );
  OR3B2S U4519 ( .I1(n5343), .B1(n5342), .B2(n5341), .O(n5349) );
  OR3B2S U4520 ( .I1(n4283), .B1(n4280), .B2(n4282), .O(n5145) );
  ND3S U4521 ( .I1(SRAM_192X32_addr[0]), .I2(SRAM_192X32_addr[1]), .I3(n4064), 
        .O(n4065) );
  AOI22S U4522 ( .A1(n5020), .A2(n5019), .B1(n5021), .B2(n3508), .O(n3643) );
  ND3S U4523 ( .I1(n5335), .I2(n5334), .I3(n5333), .O(n5337) );
  OR3B2S U4524 ( .I1(n5422), .B1(n5421), .B2(n5420), .O(n5427) );
  FA1S U4525 ( .A(n3874), .B(n3873), .CI(n3872), .CO(n3947), .S(n3950) );
  NR2 U4526 ( .I1(current_action_idx[2]), .I2(n5662), .O(n4171) );
  OR2S U4527 ( .I1(n5078), .I2(n3506), .O(n5084) );
  NR2P U4528 ( .I1(image_size_temp[0]), .I2(n3505), .O(n5755) );
  INV1S U4529 ( .I(n4938), .O(n4914) );
  INV1S U4530 ( .I(n5790), .O(n5816) );
  NR2P U4531 ( .I1(n5692), .I2(n5690), .O(n6243) );
  FA1S U4532 ( .A(n3760), .B(n3759), .CI(n3758), .CO(n3814), .S(n3831) );
  MOAI1S U4533 ( .A1(n5520), .A2(median_in[57]), .B1(n5520), .B2(n5534), .O(
        n4332) );
  FA1S U4534 ( .A(n5032), .B(n5031), .CI(n5030), .CO(n5021), .S(n5036) );
  HA1 U4535 ( .A(n6268), .B(n6267), .C(n3672), .S(n6269) );
  OA12 U4536 ( .B1(in_valid), .B2(in_valid_reg), .A1(n4209), .O(n6210) );
  MOAI1S U4537 ( .A1(n5259), .A2(median_in[8]), .B1(n5259), .B2(n5260), .O(
        n5277) );
  MOAI1S U4538 ( .A1(n5259), .A2(median_in[9]), .B1(n5259), .B2(n5264), .O(
        n4274) );
  INV1S U4539 ( .I(median_in[10]), .O(n5265) );
  INV1S U4540 ( .I(median_in[35]), .O(n5890) );
  INV1S U4541 ( .I(median_in[21]), .O(n5919) );
  OAI22S U4542 ( .A1(n5544), .A2(n5543), .B1(n5944), .B2(n5542), .O(n5554) );
  ND3S U4543 ( .I1(n5011), .I2(n5678), .I3(n5667), .O(n5055) );
  INV1S U4544 ( .I(n5095), .O(n5654) );
  FA1S U4545 ( .A(image[6]), .B(wgt_temp[5]), .CI(n5620), .CO(n5623), .S(n5622) );
  OAI12HS U4546 ( .B1(n3517), .B2(n5592), .A1(n5591), .O(n5600) );
  ND3S U4547 ( .I1(state[3]), .I2(n4068), .I3(n4067), .O(n5559) );
  FA1S U4548 ( .A(n3978), .B(n3977), .CI(n3976), .CO(mult_x_231_n48), .S(n3980) );
  ND3S U4549 ( .I1(n4462), .I2(n4461), .I3(n4460), .O(n2929) );
  ND3S U4550 ( .I1(n4436), .I2(n4435), .I3(n4434), .O(n2977) );
  ND3S U4551 ( .I1(n4080), .I2(n4168), .I3(n5557), .O(n3402) );
  ND3S U4552 ( .I1(n5936), .I2(n5206), .I3(n5205), .O(find_median_inst_max2[7]) );
  ND3S U4553 ( .I1(n4984), .I2(n4106), .I3(n4983), .O(n3000) );
  ND3S U4554 ( .I1(n4478), .I2(n4477), .I3(n4476), .O(n3121) );
  ND3S U4555 ( .I1(n4493), .I2(n4492), .I3(n4491), .O(n3115) );
  ND3S U4556 ( .I1(n4487), .I2(n4486), .I3(n4485), .O(n3109) );
  ND3S U4557 ( .I1(n4675), .I2(n4674), .I3(n4673), .O(n3026) );
  ND3S U4558 ( .I1(n4475), .I2(n4474), .I3(n4473), .O(n3059) );
  FA1S U4559 ( .A(n3970), .B(n3969), .CI(n3968), .CO(n3965), .S(N6117) );
  TIE1 U4560 ( .O(n2863) );
  OAI12HS U4561 ( .B1(n6204), .B2(avg_temp[2]), .A1(n3498), .O(n6206) );
  OAI22S U4562 ( .A1(n4582), .A2(n4617), .B1(n4581), .B2(n4617), .O(n4584) );
  OAI12HS U4563 ( .B1(n4213), .B2(avg_temp[6]), .A1(n3497), .O(n4216) );
  AOI12HS U4564 ( .B1(n3660), .B2(n4619), .A1(n5067), .O(n3658) );
  OAI12H U4565 ( .B1(n4231), .B2(n4647), .A1(n4386), .O(n5933) );
  INV1S U4566 ( .I(n4553), .O(n5725) );
  NR2 U4567 ( .I1(cal_count[4]), .I2(cal_count[5]), .O(n4004) );
  INV1S U4568 ( .I(cal_count[7]), .O(n4190) );
  ND2S U4569 ( .I1(n3488), .I2(n4190), .O(n4094) );
  NR2T U4570 ( .I1(cal_count[8]), .I2(n3984), .O(n4087) );
  INV2 U4571 ( .I(n4087), .O(n4101) );
  NR2P U4572 ( .I1(cal_count[3]), .I2(n4101), .O(n4392) );
  INV1S U4573 ( .I(n4392), .O(n4379) );
  INV1S U4574 ( .I(cal_count[0]), .O(n5692) );
  NR2 U4575 ( .I1(cal_count[2]), .I2(n6243), .O(n4090) );
  NR2 U4576 ( .I1(n4379), .I2(n4967), .O(n3661) );
  ND2S U4577 ( .I1(n3516), .I2(n3661), .O(n3520) );
  INV2 U4578 ( .I(wait_conv_out_count[1]), .O(n6070) );
  NR2P U4579 ( .I1(n6302), .I2(n6070), .O(n6069) );
  NR2 U4580 ( .I1(n6304), .I2(wait_conv_out_count[4]), .O(n3518) );
  INV1S U4581 ( .I(wait_conv_out_count[3]), .O(n3883) );
  INV2 U4582 ( .I(state[1]), .O(n4067) );
  ND2P U4583 ( .I1(n4069), .I2(state[2]), .O(n3993) );
  AOI13HS U4584 ( .B1(n6069), .B2(n3518), .B3(n3883), .A1(n3517), .O(n3519) );
  AN2 U4585 ( .I1(n3520), .I2(n3519), .O(n5695) );
  AN3B2S U4586 ( .I1(start_write_flag), .B1(SRAM_192_32_in_count[1]), .B2(
        SRAM_192_32_in_count[0]), .O(n6299) );
  ND2 U4587 ( .I1(n5692), .I2(cal_count[1]), .O(n5746) );
  NR2 U4588 ( .I1(cal_count[2]), .I2(n4945), .O(n3547) );
  INV1S U4589 ( .I(cal_count[5]), .O(n5686) );
  ND2S U4590 ( .I1(n5686), .I2(cal_count[4]), .O(n3523) );
  NR3 U4591 ( .I1(n4094), .I2(n3523), .I3(cal_count[8]), .O(n3525) );
  INV1S U4592 ( .I(n4613), .O(n5720) );
  NR2 U4593 ( .I1(cal_count[8]), .I2(cal_count[7]), .O(n4005) );
  ND3S U4594 ( .I1(n4004), .I2(n3489), .I3(n4005), .O(n4605) );
  INV1S U4595 ( .I(cal_count[8]), .O(n5656) );
  NR2 U4596 ( .I1(n5656), .I2(n3984), .O(n5748) );
  NR2F U4597 ( .I1(image_size_temp[1]), .I2(n6309), .O(n5753) );
  MOAI1 U4598 ( .A1(n5755), .A2(n4605), .B1(n5748), .B2(n3486), .O(n5723) );
  OR2 U4599 ( .I1(n5755), .I2(n5753), .O(n5766) );
  NR2 U4600 ( .I1(n4045), .I2(n4604), .O(n4610) );
  AOI13HS U4601 ( .B1(n5727), .B2(n5725), .B3(n5720), .A1(n4610), .O(n3521) );
  INV1S U4602 ( .I(n3537), .O(n3648) );
  NR2 U4603 ( .I1(n3648), .I2(state[0]), .O(n5767) );
  NR2 U4604 ( .I1(n3521), .I2(n6245), .O(n3527) );
  INV1S U4605 ( .I(n4005), .O(n3522) );
  NR3 U4606 ( .I1(cal_count[3]), .I2(n3523), .I3(n3522), .O(n4001) );
  NR2 U4607 ( .I1(cal_count[2]), .I2(n3488), .O(n3524) );
  ND3S U4608 ( .I1(n4001), .I2(n3524), .I3(n5728), .O(n4529) );
  INV1S U4609 ( .I(state[2]), .O(n4068) );
  ND3S U4610 ( .I1(state[1]), .I2(n4069), .I3(n4068), .O(n4178) );
  NR2 U4611 ( .I1(n5669), .I2(n4178), .O(n5744) );
  ND2S U4612 ( .I1(n5744), .I2(n5755), .O(n5679) );
  INV1S U4613 ( .I(n3525), .O(n3981) );
  NR2 U4614 ( .I1(cal_count[3]), .I2(n3981), .O(n4091) );
  ND3S U4615 ( .I1(cal_count[2]), .I2(n5728), .I3(n4091), .O(n4546) );
  INV1S U4616 ( .I(n4546), .O(n3526) );
  ND2S U4617 ( .I1(image_size_temp[0]), .I2(n5744), .O(n5682) );
  NR2 U4618 ( .I1(n5682), .I2(image_size_temp[1]), .O(n4545) );
  MOAI1S U4619 ( .A1(n4529), .A2(n5679), .B1(n3526), .B2(n4545), .O(n4601) );
  NR2 U4620 ( .I1(n3527), .I2(n4601), .O(n4632) );
  INV1S U4621 ( .I(n5744), .O(n3647) );
  NR2 U4622 ( .I1(n4230), .I2(n3647), .O(n3529) );
  INV1S U4623 ( .I(cal_count_5[1]), .O(n5714) );
  NR2 U4624 ( .I1(cal_count_5[2]), .I2(n5714), .O(n5994) );
  INV1S U4625 ( .I(cal_count[2]), .O(n4969) );
  NR2 U4626 ( .I1(cal_count[0]), .I2(cal_count[1]), .O(n5729) );
  OAI12HS U4627 ( .B1(n4969), .B2(n5729), .A1(n4392), .O(n3528) );
  NR2 U4628 ( .I1(n4553), .I2(n4608), .O(n5721) );
  AO12S U4629 ( .B1(n5766), .B2(n5729), .A1(n5721), .O(n3530) );
  ND3S U4630 ( .I1(n5767), .I2(n4101), .I3(n3530), .O(n3531) );
  XOR2HS U4631 ( .I1(rd_addr[7]), .I2(action_reg_0__1_), .O(n3536) );
  INV1S U4632 ( .I(action_reg_0__0_), .O(n3534) );
  INV1S U4633 ( .I(rd_addr[6]), .O(n3533) );
  NR2 U4634 ( .I1(n3534), .I2(n3533), .O(n3535) );
  XOR2HS U4635 ( .I1(n3536), .I2(n3535), .O(n3667) );
  NR2 U4636 ( .I1(n4230), .I2(n3549), .O(n3649) );
  AN2 U4637 ( .I1(state[0]), .I2(flip_flag), .O(n4539) );
  ND2P U4638 ( .I1(n3537), .I2(n4539), .O(n4082) );
  NR2 U4639 ( .I1(n4101), .I2(n5745), .O(n4527) );
  ND2S U4640 ( .I1(n5728), .I2(n4527), .O(n3551) );
  INV1S U4641 ( .I(n3551), .O(n4541) );
  ND3S U4642 ( .I1(n3649), .I2(n4542), .I3(n4541), .O(n3631) );
  INV1S U4643 ( .I(n3631), .O(n3539) );
  ND3S U4644 ( .I1(n4392), .I2(cal_count[2]), .I3(n5728), .O(n4540) );
  INV1S U4645 ( .I(n5755), .O(n5751) );
  ND2S U4646 ( .I1(n3660), .I2(n4539), .O(n3554) );
  NR2 U4647 ( .I1(n4540), .I2(n3554), .O(n3538) );
  ND3S U4648 ( .I1(n4087), .I2(n3547), .I3(n5728), .O(n4582) );
  NR2 U4649 ( .I1(n4582), .I2(n3554), .O(n3632) );
  OR2 U4650 ( .I1(n3538), .I2(n3632), .O(n3638) );
  INV1S U4651 ( .I(n6299), .O(n4787) );
  NR2 U4652 ( .I1(n5610), .I2(n4787), .O(n4786) );
  AN2 U4653 ( .I1(n4786), .I2(n5095), .O(n3637) );
  INV1S U4654 ( .I(n3637), .O(n3630) );
  INV1S U4655 ( .I(SRAM_192X32_addr[7]), .O(n3581) );
  INV1S U4656 ( .I(n3561), .O(n3541) );
  INV1S U4657 ( .I(n3657), .O(n3540) );
  ND2S U4658 ( .I1(n3541), .I2(n3577), .O(n3663) );
  AN2 U4659 ( .I1(n3663), .I2(n5984), .O(n3622) );
  MOAI1S U4660 ( .A1(n3630), .A2(n3581), .B1(n3622), .B2(wb_addr[7]), .O(n3542) );
  OR2 U4661 ( .I1(n3637), .I2(n3628), .O(n5080) );
  INV1S U4662 ( .I(n5745), .O(n4376) );
  ND3S U4663 ( .I1(n4087), .I2(n5727), .I3(n4376), .O(n4581) );
  NR2 U4664 ( .I1(n4581), .I2(n4542), .O(n4550) );
  INV1S U4665 ( .I(n4550), .O(n3543) );
  OR2S U4666 ( .I1(n3543), .I2(n3662), .O(n3546) );
  NR2 U4667 ( .I1(n4581), .I2(n4082), .O(n4569) );
  OAI12HS U4668 ( .B1(n4582), .B2(n4542), .A1(n3550), .O(n4549) );
  ND2S U4669 ( .I1(n3660), .I2(n4549), .O(n3545) );
  INV1S U4670 ( .I(cal_count_5[0]), .O(n4986) );
  ND2S U4671 ( .I1(n3561), .I2(n5985), .O(n3544) );
  ND3S U4672 ( .I1(n3546), .I2(n3545), .I3(n3544), .O(n3613) );
  INV1S U4673 ( .I(n3982), .O(n3548) );
  ND2S U4674 ( .I1(n4087), .I2(n3548), .O(n4563) );
  NR2 U4675 ( .I1(cal_count_5[2]), .I2(n5710), .O(n5743) );
  NR2 U4676 ( .I1(n4101), .I2(n4387), .O(n3570) );
  OR2S U4677 ( .I1(n6243), .I2(n3570), .O(n4570) );
  NR2 U4678 ( .I1(n4553), .I2(n3549), .O(n3665) );
  AOI22S U4679 ( .A1(n5743), .A2(n3663), .B1(n4570), .B2(n3665), .O(n3553) );
  NR2 U4680 ( .I1(n4542), .I2(n3551), .O(n4564) );
  OAI12HS U4681 ( .B1(n4569), .B2(n4564), .A1(n3649), .O(n3552) );
  OAI112HS U4682 ( .C1(n3554), .C2(n4563), .A1(n3553), .B1(n3552), .O(n3555)
         );
  NR2 U4683 ( .I1(n3613), .I2(n3555), .O(n3621) );
  INV1S U4684 ( .I(n3660), .O(n3573) );
  INV1S U4685 ( .I(n5750), .O(n3556) );
  NR2 U4686 ( .I1(n4969), .I2(n4945), .O(n4003) );
  AOI13HS U4687 ( .B1(cal_count[5]), .B2(n3556), .B3(n5688), .A1(cal_count[8]), 
        .O(n3568) );
  NR2 U4688 ( .I1(n4003), .I2(n4101), .O(n4618) );
  INV1S U4689 ( .I(n4618), .O(n3557) );
  INV1S U4690 ( .I(n3567), .O(n3558) );
  NR2 U4691 ( .I1(n3573), .I2(n4585), .O(n3601) );
  ND2S U4692 ( .I1(cal_count[2]), .I2(n5727), .O(n4381) );
  NR2 U4693 ( .I1(n4379), .I2(n4381), .O(n4095) );
  INV1S U4694 ( .I(n4095), .O(n3559) );
  OAI12HS U4695 ( .B1(n4540), .B2(n4542), .A1(n3559), .O(n4556) );
  ND2S U4696 ( .I1(n4556), .I2(n3660), .O(n3564) );
  NR2 U4697 ( .I1(cal_count_5[0]), .I2(cal_count_5[1]), .O(n6028) );
  INV1S U4698 ( .I(cal_count_5[2]), .O(n6024) );
  NR2 U4699 ( .I1(n5746), .I2(n4527), .O(n5758) );
  INV1S U4700 ( .I(n3662), .O(n3560) );
  AOI22S U4701 ( .A1(n6016), .A2(n3561), .B1(n4555), .B2(n3560), .O(n3563) );
  INV1S U4702 ( .I(n5729), .O(n4621) );
  ND2S U4703 ( .I1(n4554), .I2(n3665), .O(n3562) );
  ND3S U4704 ( .I1(n3564), .I2(n3563), .I3(n3562), .O(n3617) );
  NR2 U4705 ( .I1(n3601), .I2(n3617), .O(n3579) );
  ND3S U4706 ( .I1(cal_count[5]), .I2(n3489), .I3(cal_count[7]), .O(n4187) );
  NR2 U4707 ( .I1(n4187), .I2(n4945), .O(n3565) );
  ND3S U4708 ( .I1(n3565), .I2(cal_count[4]), .I3(n4967), .O(n3566) );
  ND2S U4709 ( .I1(n5656), .I2(n3566), .O(n4606) );
  NR2 U4710 ( .I1(n4618), .I2(n4606), .O(n3659) );
  MOAI1S U4711 ( .A1(n3568), .A2(n3567), .B1(n5727), .B2(n3659), .O(n3569) );
  INV1S U4712 ( .I(n6243), .O(n4943) );
  INV1S U4713 ( .I(n3577), .O(n3571) );
  MOAI1S U4714 ( .A1(n3662), .A2(n4943), .B1(n3571), .B2(n6016), .O(n3572) );
  AOI12HS U4715 ( .B1(n4532), .B2(n3660), .A1(n3572), .O(n3578) );
  NR2 U4716 ( .I1(n4542), .I2(n4563), .O(n4534) );
  ND2S U4717 ( .I1(n4095), .I2(n4082), .O(n4535) );
  NR2 U4718 ( .I1(n3573), .I2(n4535), .O(n3574) );
  NR2 U4719 ( .I1(n3623), .I2(n3574), .O(n3618) );
  INV1S U4720 ( .I(n5985), .O(n3576) );
  ND2S U4721 ( .I1(n3660), .I2(n4550), .O(n3575) );
  AN3 U4722 ( .I1(n3578), .I2(n3618), .I3(n3507), .O(n3609) );
  ND3 U4723 ( .I1(n3621), .I2(n3579), .I3(n3609), .O(n3641) );
  INV1S U4724 ( .I(n5610), .O(n4209) );
  INV1S U4725 ( .I(RGB_count[1]), .O(n3675) );
  INV1S U4726 ( .I(RGB_count[0]), .O(n3898) );
  NR2 U4727 ( .I1(n3675), .I2(n3898), .O(n3676) );
  NR2 U4728 ( .I1(n3676), .I2(n4787), .O(n4788) );
  NR2 U4729 ( .I1(n4209), .I2(n3580), .O(n3639) );
  INV1S U4730 ( .I(n3639), .O(n3590) );
  INV1S U4731 ( .I(n3622), .O(n3597) );
  MOAI1S U4732 ( .A1(n3590), .A2(n3581), .B1(n3622), .B2(action_reg_0__1_), 
        .O(n3582) );
  XOR2HS U4733 ( .I1(n5080), .I2(n3583), .O(n3584) );
  XOR2HS U4734 ( .I1(n3585), .I2(n3584), .O(n3644) );
  XOR2HS U4735 ( .I1(action_reg_0__0_), .I2(rd_addr[6]), .O(n5026) );
  ND2S U4736 ( .I1(n3622), .I2(action_reg_0__0_), .O(n3587) );
  ND2S U4737 ( .I1(n3639), .I2(SRAM_192X32_addr[6]), .O(n3586) );
  XOR2HS U4738 ( .I1(n5080), .I2(n3589), .O(n5020) );
  ND2S U4739 ( .I1(n3622), .I2(wb_addr[6]), .O(n3591) );
  OAI112HS U4740 ( .C1(n3630), .C2(n6303), .A1(n3591), .B1(n3590), .O(n3592)
         );
  INV1S U4741 ( .I(wb_addr[5]), .O(n3593) );
  MOAI1S U4742 ( .A1(n3597), .A2(n3593), .B1(n3637), .B2(SRAM_192X32_addr[5]), 
        .O(n3594) );
  XOR2HS U4743 ( .I1(n5080), .I2(n3596), .O(n5031) );
  INV1S U4744 ( .I(wb_addr[4]), .O(n5041) );
  MOAI1S U4745 ( .A1(n3597), .A2(n5041), .B1(n3637), .B2(SRAM_192X32_addr[4]), 
        .O(n3598) );
  XOR2HS U4746 ( .I1(n5080), .I2(n3600), .O(n5090) );
  INV1S U4747 ( .I(n3601), .O(n3604) );
  ND2S U4748 ( .I1(n3622), .I2(wb_addr[3]), .O(n3603) );
  ND2S U4749 ( .I1(n3637), .I2(SRAM_192X32_addr[3]), .O(n3602) );
  XOR2HS U4750 ( .I1(n5080), .I2(n3607), .O(n5044) );
  AOI22S U4751 ( .A1(n3637), .A2(SRAM_192X32_addr[2]), .B1(n3622), .B2(
        wb_addr[2]), .O(n3608) );
  ND2S U4752 ( .I1(n3609), .I2(n3608), .O(n3610) );
  AO12S U4753 ( .B1(n3639), .B2(SRAM_192X32_addr[2]), .A1(n3637), .O(n3611) );
  XOR2HS U4754 ( .I1(n5080), .I2(n3612), .O(n5057) );
  INV1S U4755 ( .I(n3613), .O(n3615) );
  AOI22S U4756 ( .A1(n3637), .A2(SRAM_192X32_addr[1]), .B1(n3622), .B2(
        wb_addr[1]), .O(n3614) );
  ND2S U4757 ( .I1(n3615), .I2(n3614), .O(n3616) );
  NR2 U4758 ( .I1(n3617), .I2(n3616), .O(n3619) );
  ND2S U4759 ( .I1(n3619), .I2(n3618), .O(n3620) );
  ND2S U4760 ( .I1(n3622), .I2(wb_addr[0]), .O(n3625) );
  ND2S U4761 ( .I1(n3637), .I2(SRAM_192X32_addr[0]), .O(n3624) );
  AN4B1S U4762 ( .I1(n3507), .I2(n3625), .I3(n3624), .B1(n3623), .O(n3626) );
  ND2S U4763 ( .I1(n3621), .I2(n3626), .O(n3627) );
  NR2 U4764 ( .I1(n5080), .I2(n5079), .O(n3636) );
  ND2S U4765 ( .I1(n3639), .I2(SRAM_192X32_addr[0]), .O(n3629) );
  ND3S U4766 ( .I1(n3631), .I2(n3630), .I3(n3629), .O(n3633) );
  OR2S U4767 ( .I1(n3633), .I2(n3632), .O(n3634) );
  AO12 U4768 ( .B1(N1043), .B2(n3641), .A1(n3634), .O(n3635) );
  XNR2HS U4769 ( .I1(n5080), .I2(n3635), .O(n5082) );
  MOAI1 U4770 ( .A1(n3636), .A2(n5082), .B1(n5079), .B2(n5080), .O(n5070) );
  AO112S U4771 ( .C1(n3639), .C2(SRAM_192X32_addr[1]), .A1(n3638), .B1(n3637), 
        .O(n3640) );
  XOR2HS U4772 ( .I1(n5080), .I2(n3642), .O(n5069) );
  XNR2HS U4773 ( .I1(n3644), .I2(n3643), .O(n3655) );
  INV1S U4774 ( .I(n6028), .O(n3645) );
  ND3S U4775 ( .I1(n3646), .I2(n5744), .I3(n5766), .O(n4597) );
  NR2 U4776 ( .I1(action_idx[3]), .I2(action_idx[2]), .O(n5580) );
  INV1S U4777 ( .I(n5580), .O(n5585) );
  NR2 U4778 ( .I1(action_idx[0]), .I2(n5585), .O(n3991) );
  INV1S U4779 ( .I(action_idx[1]), .O(n5576) );
  ND3S U4780 ( .I1(n3537), .I2(n6309), .I3(n4608), .O(n3651) );
  INV1S U4781 ( .I(n3649), .O(n3650) );
  OAI22S U4782 ( .A1(n6299), .A2(n3651), .B1(n4554), .B2(n3650), .O(n3652) );
  MOAI1S U4783 ( .A1(n6299), .A2(n3653), .B1(n6301), .B2(n3652), .O(n3654) );
  NR3 U4784 ( .I1(n5654), .I2(n4788), .I3(n3654), .O(n5093) );
  INV1S U4785 ( .I(n5093), .O(n5098) );
  AN2B1S U4786 ( .I1(n3657), .B1(n3656), .O(n5067) );
  NR2 U4787 ( .I1(n4376), .I2(n4101), .O(n4089) );
  MOAI1S U4788 ( .A1(n4003), .A2(n4378), .B1(n5729), .B2(n4089), .O(n4619) );
  NR2 U4789 ( .I1(n5093), .I2(n3658), .O(n5024) );
  AOI22S U4790 ( .A1(n5093), .A2(SRAM_192X32_addr[7]), .B1(n5024), .B2(
        action_reg_0__1_), .O(n3669) );
  MOAI1S U4791 ( .A1(n3662), .A2(n3661), .B1(n3660), .B2(n3659), .O(n3664) );
  INV1S U4792 ( .I(n5713), .O(n6015) );
  INV1S U4793 ( .I(avg_temp[9]), .O(n4210) );
  AN2S U4794 ( .I1(n5610), .I2(avg_temp[8]), .O(n6268) );
  AN2S U4795 ( .I1(n5610), .I2(avg_temp[7]), .O(n6271) );
  MOAI1S U4796 ( .A1(n3672), .A2(n3671), .B1(n3672), .B2(n3671), .O(n3673) );
  MOAI1 U4797 ( .A1(n3493), .A2(n4210), .B1(n3493), .B2(n3673), .O(n2615) );
  NR2 U4798 ( .I1(n5134), .I2(n5626), .O(n5624) );
  INV1S U4799 ( .I(n5624), .O(n3677) );
  INV1S U4800 ( .I(median_in[49]), .O(n5526) );
  INV1S U4801 ( .I(n6071), .O(n5106) );
  NR2P U4802 ( .I1(wait_conv_out_count[4]), .I2(n3883), .O(n3684) );
  ND3S U4803 ( .I1(n5106), .I2(N6291), .I3(n3684), .O(n3767) );
  NR2 U4804 ( .I1(n6304), .I2(n6070), .O(n6090) );
  ND3S U4805 ( .I1(n6090), .I2(n3684), .I3(n6302), .O(n3692) );
  INV1S U4806 ( .I(median_in[33]), .O(n5177) );
  OAI22S U4807 ( .A1(n5526), .A2(n3767), .B1(n3692), .B2(n5177), .O(n3683) );
  INV1S U4808 ( .I(median_in[17]), .O(n5264) );
  NR2 U4809 ( .I1(N6291), .I2(wait_conv_out_count[3]), .O(n61150) );
  ND2S U4810 ( .I1(n61150), .I2(wait_conv_out_count[4]), .O(n6114) );
  NR2 U4811 ( .I1(n3679), .I2(n6114), .O(n3680) );
  BUF2 U4812 ( .I(n3680), .O(n3799) );
  MOAI1S U4813 ( .A1(n5264), .A2(n3768), .B1(n3799), .B2(median_in[1]), .O(
        n3682) );
  INV1S U4814 ( .I(median_in[57]), .O(n5525) );
  INV1S U4815 ( .I(n6069), .O(n4957) );
  NR2 U4816 ( .I1(N6291), .I2(n4957), .O(n4961) );
  ND2S U4817 ( .I1(n4961), .I2(n3684), .O(n3691) );
  INV1S U4818 ( .I(median_in[65]), .O(n5534) );
  NR2 U4819 ( .I1(N6291), .I2(n6070), .O(n6093) );
  OAI22S U4820 ( .A1(n5525), .A2(n3691), .B1(n5534), .B2(n3769), .O(n3681) );
  NR3 U4821 ( .I1(n3683), .I2(n3682), .I3(n3681), .O(n3689) );
  NR2 U4822 ( .I1(n6304), .I2(wait_conv_out_count[1]), .O(n6107) );
  NR2 U4823 ( .I1(n6083), .I2(n4957), .O(n4948) );
  INV1S U4824 ( .I(wait_conv_out_count[4]), .O(n5105) );
  ND2P U4825 ( .I1(n4948), .I2(n5105), .O(n4951) );
  INV1S U4826 ( .I(n4951), .O(n3773) );
  AOI22S U4827 ( .A1(n3789), .A2(median_in[41]), .B1(n3773), .B2(median_in[25]), .O(n3688) );
  NR2 U4828 ( .I1(n3685), .I2(n6114), .O(n3686) );
  ND3S U4829 ( .I1(n3689), .I2(n3688), .I3(n3687), .O(n3690) );
  INV1S U4830 ( .I(n3690), .O(n3836) );
  INV2 U4831 ( .I(n3769), .O(n3795) );
  INV2 U4832 ( .I(n3691), .O(n3699) );
  AOI22S U4833 ( .A1(n3795), .A2(template_reg[69]), .B1(n3699), .B2(
        template_reg[61]), .O(n3695) );
  INV2 U4834 ( .I(n3692), .O(n3797) );
  INV2 U4835 ( .I(n3767), .O(n3796) );
  AOI22S U4836 ( .A1(n3797), .A2(template_reg[37]), .B1(n3796), .B2(
        template_reg[53]), .O(n3694) );
  INV2 U4837 ( .I(n3768), .O(n3798) );
  AOI22S U4838 ( .A1(n3799), .A2(template_reg[5]), .B1(n3798), .B2(
        template_reg[21]), .O(n3693) );
  ND3S U4839 ( .I1(n3695), .I2(n3694), .I3(n3693), .O(n3698) );
  INV1S U4840 ( .I(template_reg[29]), .O(n3696) );
  MOAI1S U4841 ( .A1(n4951), .A2(n3696), .B1(n3789), .B2(template_reg[45]), 
        .O(n3697) );
  NR2 U4842 ( .I1(n3836), .I2(n3502), .O(n3809) );
  INV1S U4843 ( .I(median_in[51]), .O(n5893) );
  MOAI1S U4844 ( .A1(n5893), .A2(n3767), .B1(n3797), .B2(median_in[35]), .O(
        n3702) );
  INV1S U4845 ( .I(median_in[19]), .O(n5268) );
  MOAI1S U4846 ( .A1(n5268), .A2(n3768), .B1(n3799), .B2(median_in[3]), .O(
        n3701) );
  INV1S U4847 ( .I(median_in[67]), .O(n5894) );
  MOAI1S U4848 ( .A1(n5894), .A2(n3769), .B1(n3699), .B2(median_in[59]), .O(
        n3700) );
  NR3 U4849 ( .I1(n3702), .I2(n3701), .I3(n3700), .O(n3705) );
  AOI22S U4850 ( .A1(n3789), .A2(median_in[43]), .B1(n3773), .B2(median_in[27]), .O(n3704) );
  AOI22S U4851 ( .A1(template_reg[67]), .A2(n3795), .B1(n3699), .B2(
        template_reg[59]), .O(n3708) );
  AOI22S U4852 ( .A1(n3797), .A2(template_reg[35]), .B1(n3796), .B2(
        template_reg[51]), .O(n3707) );
  AOI22S U4853 ( .A1(n3799), .A2(template_reg[3]), .B1(n3798), .B2(
        template_reg[19]), .O(n3706) );
  ND3S U4854 ( .I1(n3708), .I2(n3707), .I3(n3706), .O(n3711) );
  INV1S U4855 ( .I(template_reg[27]), .O(n3709) );
  MOAI1S U4856 ( .A1(n4951), .A2(n3709), .B1(template_reg[43]), .B2(n3789), 
        .O(n3710) );
  NR2 U4857 ( .I1(n3511), .I2(n3496), .O(n3808) );
  AOI22S U4858 ( .A1(median_in[66]), .A2(n3795), .B1(n3699), .B2(median_in[58]), .O(n3714) );
  AOI22S U4859 ( .A1(n3797), .A2(median_in[34]), .B1(n3796), .B2(median_in[50]), .O(n3713) );
  AOI22S U4860 ( .A1(n3799), .A2(median_in[2]), .B1(n3798), .B2(median_in[18]), 
        .O(n3712) );
  ND3S U4861 ( .I1(n3714), .I2(n3713), .I3(n3712), .O(n3716) );
  MOAI1S U4862 ( .A1(n4951), .A2(n6318), .B1(median_in[42]), .B2(n3789), .O(
        n3715) );
  AOI22S U4863 ( .A1(template_reg[68]), .A2(n3795), .B1(n3699), .B2(
        template_reg[60]), .O(n3719) );
  AOI22S U4864 ( .A1(n3797), .A2(template_reg[36]), .B1(n3796), .B2(
        template_reg[52]), .O(n3718) );
  AOI22S U4865 ( .A1(n3799), .A2(template_reg[4]), .B1(n3798), .B2(
        template_reg[20]), .O(n3717) );
  ND3S U4866 ( .I1(n3719), .I2(n3718), .I3(n3717), .O(n3722) );
  INV1S U4867 ( .I(template_reg[28]), .O(n3720) );
  MOAI1S U4868 ( .A1(n4951), .A2(n3720), .B1(template_reg[44]), .B2(n3789), 
        .O(n3721) );
  NR2 U4869 ( .I1(n3512), .I2(n3503), .O(n3807) );
  NR2 U4870 ( .I1(n3836), .I2(n3503), .O(n3760) );
  NR2 U4871 ( .I1(n3512), .I2(n3496), .O(n3759) );
  INV1S U4872 ( .I(median_in[52]), .O(n5904) );
  MOAI1S U4873 ( .A1(n5904), .A2(n3767), .B1(n3797), .B2(median_in[36]), .O(
        n3725) );
  INV1S U4874 ( .I(median_in[20]), .O(n5909) );
  MOAI1S U4875 ( .A1(n5909), .A2(n3768), .B1(n3799), .B2(median_in[4]), .O(
        n3724) );
  INV1S U4876 ( .I(median_in[68]), .O(n5532) );
  MOAI1S U4877 ( .A1(n5532), .A2(n3769), .B1(n3699), .B2(median_in[60]), .O(
        n3723) );
  NR3 U4878 ( .I1(n3725), .I2(n3724), .I3(n3723), .O(n3728) );
  AOI22S U4879 ( .A1(n3789), .A2(median_in[44]), .B1(n3773), .B2(median_in[28]), .O(n3727) );
  ND3S U4880 ( .I1(n3728), .I2(n3727), .I3(n3726), .O(n3729) );
  INV1S U4881 ( .I(n3729), .O(n3854) );
  AOI22S U4882 ( .A1(template_reg[65]), .A2(n3795), .B1(n3699), .B2(
        template_reg[57]), .O(n3732) );
  AOI22S U4883 ( .A1(n3797), .A2(template_reg[33]), .B1(n3796), .B2(
        template_reg[49]), .O(n3731) );
  AOI22S U4884 ( .A1(n3799), .A2(template_reg[1]), .B1(n3798), .B2(
        template_reg[17]), .O(n3730) );
  ND3S U4885 ( .I1(n3732), .I2(n3731), .I3(n3730), .O(n3735) );
  INV1S U4886 ( .I(template_reg[25]), .O(n3733) );
  MOAI1S U4887 ( .A1(n4951), .A2(n3733), .B1(template_reg[41]), .B2(n3789), 
        .O(n3734) );
  NR2 U4888 ( .I1(n3854), .I2(n3501), .O(n3782) );
  AOI22S U4889 ( .A1(n3795), .A2(median_in[69]), .B1(n3699), .B2(median_in[61]), .O(n3738) );
  AOI22S U4890 ( .A1(n3797), .A2(median_in[37]), .B1(median_in[53]), .B2(n3796), .O(n3737) );
  AOI22S U4891 ( .A1(n3799), .A2(median_in[5]), .B1(n3798), .B2(median_in[21]), 
        .O(n3736) );
  ND3S U4892 ( .I1(n3738), .I2(n3737), .I3(n3736), .O(n3740) );
  INV1S U4893 ( .I(median_in[29]), .O(n5179) );
  INV1S U4894 ( .I(median_in[45]), .O(n5184) );
  OAI22S U4895 ( .A1(n5179), .A2(n4951), .B1(n5184), .B2(n3803), .O(n3739) );
  AOI22S U4896 ( .A1(template_reg[64]), .A2(n3795), .B1(n3699), .B2(
        template_reg[56]), .O(n3743) );
  AOI22S U4897 ( .A1(n3797), .A2(template_reg[32]), .B1(n3796), .B2(
        template_reg[48]), .O(n3742) );
  AOI22S U4898 ( .A1(n3799), .A2(template_reg[0]), .B1(n3798), .B2(
        template_reg[16]), .O(n3741) );
  ND3S U4899 ( .I1(n3743), .I2(n3742), .I3(n3741), .O(n3746) );
  INV1S U4900 ( .I(template_reg[24]), .O(n3744) );
  MOAI1S U4901 ( .A1(n4951), .A2(n3744), .B1(template_reg[40]), .B2(n3789), 
        .O(n3745) );
  NR2 U4902 ( .I1(n3510), .I2(n3494), .O(n3781) );
  AOI22S U4903 ( .A1(median_in[64]), .A2(n3795), .B1(n3699), .B2(median_in[56]), .O(n3749) );
  AOI22S U4904 ( .A1(n3797), .A2(median_in[32]), .B1(n3796), .B2(median_in[48]), .O(n3748) );
  AOI22S U4905 ( .A1(n3799), .A2(median_in[0]), .B1(n3798), .B2(median_in[16]), 
        .O(n3747) );
  ND3S U4906 ( .I1(n3749), .I2(n3748), .I3(n3747), .O(n3751) );
  INV1S U4907 ( .I(median_in[24]), .O(n5176) );
  INV1S U4908 ( .I(median_in[40]), .O(n5175) );
  OAI22S U4909 ( .A1(n5176), .A2(n4951), .B1(n3803), .B2(n5175), .O(n3750) );
  NR2 U4910 ( .I1(n3515), .I2(n3503), .O(n3818) );
  AOI22S U4911 ( .A1(template_reg[66]), .A2(n3795), .B1(n3699), .B2(
        template_reg[58]), .O(n3754) );
  AOI22S U4912 ( .A1(n3797), .A2(template_reg[34]), .B1(n3796), .B2(
        template_reg[50]), .O(n3753) );
  AOI22S U4913 ( .A1(n3799), .A2(template_reg[2]), .B1(n3798), .B2(
        template_reg[18]), .O(n3752) );
  ND3S U4914 ( .I1(n3754), .I2(n3753), .I3(n3752), .O(n3757) );
  INV1S U4915 ( .I(template_reg[26]), .O(n3755) );
  MOAI1S U4916 ( .A1(n4951), .A2(n3755), .B1(template_reg[42]), .B2(n3789), 
        .O(n3756) );
  NR2 U4917 ( .I1(n3512), .I2(n3499), .O(n3817) );
  NR2 U4918 ( .I1(n3512), .I2(n3501), .O(n3822) );
  NR2 U4919 ( .I1(n3511), .I2(n3494), .O(n3821) );
  NR2 U4920 ( .I1(n3515), .I2(n3502), .O(n3780) );
  NR2 U4921 ( .I1(n3511), .I2(n3499), .O(n3779) );
  NR2 U4922 ( .I1(n3511), .I2(n3501), .O(n3820) );
  NR2 U4923 ( .I1(n3854), .I2(n3494), .O(n3819) );
  NR2 U4924 ( .I1(n3511), .I2(n3503), .O(n3862) );
  AOI22S U4925 ( .A1(n3795), .A2(template_reg[70]), .B1(n3699), .B2(
        template_reg[62]), .O(n3763) );
  AOI22S U4926 ( .A1(n3797), .A2(template_reg[38]), .B1(n3796), .B2(
        template_reg[54]), .O(n3762) );
  AOI22S U4927 ( .A1(n3799), .A2(template_reg[6]), .B1(n3798), .B2(
        template_reg[22]), .O(n3761) );
  INV1S U4928 ( .I(template_reg[30]), .O(n3764) );
  MOAI1S U4929 ( .A1(n4951), .A2(n3764), .B1(n3789), .B2(template_reg[46]), 
        .O(n3765) );
  NR2 U4930 ( .I1(n3836), .I2(n3500), .O(n3861) );
  NR2 U4931 ( .I1(n3854), .I2(n3496), .O(n3860) );
  NR2 U4932 ( .I1(n3510), .I2(n3501), .O(n3794) );
  INV1S U4933 ( .I(median_in[54]), .O(n5926) );
  INV1S U4934 ( .I(median_in[22]), .O(n5271) );
  INV1S U4935 ( .I(median_in[70]), .O(n5927) );
  MOAI1S U4936 ( .A1(n5927), .A2(n3769), .B1(n3699), .B2(median_in[62]), .O(
        n3770) );
  NR3 U4937 ( .I1(n3772), .I2(n3771), .I3(n3770), .O(n3776) );
  AOI22S U4938 ( .A1(n3789), .A2(median_in[46]), .B1(n3773), .B2(median_in[30]), .O(n3775) );
  ND3S U4939 ( .I1(n3776), .I2(n3775), .I3(n3774), .O(n3777) );
  INV1S U4940 ( .I(n3777), .O(n3910) );
  NR2 U4941 ( .I1(n3910), .I2(n3494), .O(n3793) );
  FA1 U4942 ( .A(n3780), .B(n3779), .CI(n3778), .CO(n3811), .S(n3832) );
  NR2 U4943 ( .I1(n3515), .I2(n3500), .O(n3785) );
  NR2 U4944 ( .I1(n3854), .I2(n3499), .O(n3784) );
  HA1 U4945 ( .A(n3782), .B(n3781), .C(n3783), .S(n3758) );
  FA1S U4946 ( .A(n3785), .B(n3784), .CI(n3783), .CO(n3952), .S(n3810) );
  AOI22S U4947 ( .A1(n3795), .A2(template_reg[71]), .B1(n3699), .B2(
        template_reg[63]), .O(n3788) );
  AOI22S U4948 ( .A1(n3797), .A2(template_reg[39]), .B1(n3796), .B2(
        template_reg[55]), .O(n3787) );
  AOI22S U4949 ( .A1(n3799), .A2(template_reg[7]), .B1(n3798), .B2(
        template_reg[23]), .O(n3786) );
  INV1S U4950 ( .I(template_reg[31]), .O(n3790) );
  MOAI1S U4951 ( .A1(n4951), .A2(n3790), .B1(n3789), .B2(template_reg[47]), 
        .O(n3791) );
  NR2 U4952 ( .I1(n3515), .I2(n3495), .O(n3868) );
  NR2 U4953 ( .I1(n3510), .I2(n3499), .O(n3867) );
  NR2 U4954 ( .I1(n3512), .I2(n3502), .O(n3874) );
  NR2 U4955 ( .I1(n3910), .I2(n3501), .O(n3838) );
  AOI22S U4956 ( .A1(n3795), .A2(median_in[71]), .B1(n3699), .B2(median_in[63]), .O(n3802) );
  AOI22S U4957 ( .A1(n3797), .A2(median_in[39]), .B1(n3796), .B2(median_in[55]), .O(n3801) );
  AOI22S U4958 ( .A1(n3799), .A2(median_in[7]), .B1(n3798), .B2(median_in[23]), 
        .O(n3800) );
  INV1S U4959 ( .I(median_in[31]), .O(n5206) );
  INV1S U4960 ( .I(median_in[47]), .O(n5205) );
  OAI22S U4961 ( .A1(n5206), .A2(n4951), .B1(n5205), .B2(n3803), .O(n3804) );
  NR2 U4962 ( .I1(n3509), .I2(n3494), .O(n3837) );
  FA1S U4963 ( .A(n3812), .B(n3811), .CI(n3810), .CO(n3954), .S(n3961) );
  FA1 U4964 ( .A(n3815), .B(n3814), .CI(n3813), .CO(n3958), .S(n3960) );
  NR2 U4965 ( .I1(n3836), .I2(n3496), .O(n3830) );
  NR2 U4966 ( .I1(n3515), .I2(n3496), .O(n3825) );
  NR2 U4967 ( .I1(n3836), .I2(n3499), .O(n3824) );
  NR2 U4968 ( .I1(n3515), .I2(n3499), .O(n3827) );
  NR2 U4969 ( .I1(n3836), .I2(n3501), .O(n3826) );
  FA1 U4970 ( .A(n3825), .B(n3824), .CI(n3823), .CO(n3828), .S(n3966) );
  NR2 U4971 ( .I1(n3512), .I2(n3494), .O(n3970) );
  NR2 U4972 ( .I1(n3836), .I2(n3494), .O(n3972) );
  NR2 U4973 ( .I1(n3515), .I2(n3501), .O(n3971) );
  HA1 U4974 ( .A(n3827), .B(n3826), .C(n3823), .S(n3968) );
  INV1S U4975 ( .I(n3908), .O(n3835) );
  FA1 U4976 ( .A(n3833), .B(n3832), .CI(n3831), .CO(n3813), .S(n3906) );
  NR2P U4977 ( .I1(n3907), .I2(n3906), .O(n3834) );
  NR2 U4978 ( .I1(n3854), .I2(n3502), .O(n3847) );
  NR2 U4979 ( .I1(n3836), .I2(n3495), .O(n3865) );
  NR2 U4980 ( .I1(n3511), .I2(n3502), .O(n3864) );
  NR2 U4981 ( .I1(n3512), .I2(n3500), .O(n3863) );
  NR2 U4982 ( .I1(n3854), .I2(n3503), .O(n3871) );
  NR2 U4983 ( .I1(n3510), .I2(n3496), .O(n3870) );
  HA1 U4984 ( .A(n3838), .B(n3837), .C(n3869), .S(n3873) );
  NR2 U4985 ( .I1(n3512), .I2(n3495), .O(n3844) );
  NR2 U4986 ( .I1(n3509), .I2(n3499), .O(n3843) );
  NR2 U4987 ( .I1(n3910), .I2(n3499), .O(n3859) );
  NR2 U4988 ( .I1(n3509), .I2(n3501), .O(n3858) );
  NR2 U4989 ( .I1(n3511), .I2(n3495), .O(n3853) );
  NR2 U4990 ( .I1(n3509), .I2(n3496), .O(n3852) );
  NR2 U4991 ( .I1(n3854), .I2(n3500), .O(n3851) );
  NR2 U4992 ( .I1(n3510), .I2(n3502), .O(n3850) );
  NR2 U4993 ( .I1(n3910), .I2(n3503), .O(n3849) );
  NR2 U4994 ( .I1(n3510), .I2(n3503), .O(n3841) );
  NR2 U4995 ( .I1(n3511), .I2(n3500), .O(n3840) );
  NR2 U4996 ( .I1(n3910), .I2(n3496), .O(n3839) );
  FA1S U4997 ( .A(n3841), .B(n3840), .CI(n3839), .CO(n3848), .S(n3877) );
  FA1S U4998 ( .A(n3844), .B(n3843), .CI(n3842), .CO(n3857), .S(n3876) );
  FA1S U4999 ( .A(n3847), .B(n3846), .CI(n3845), .CO(n3880), .S(n3875) );
  FA1S U5000 ( .A(n3850), .B(n3849), .CI(n3848), .CO(n3928), .S(n3855) );
  NR2 U5001 ( .I1(n3510), .I2(n3500), .O(n3922) );
  FA1S U5002 ( .A(n3853), .B(n3852), .CI(n3851), .CO(n3921), .S(n3856) );
  NR2 U5003 ( .I1(n3854), .I2(n3495), .O(n3916) );
  NR2 U5004 ( .I1(n3509), .I2(n3503), .O(n3915) );
  NR2 U5005 ( .I1(n3910), .I2(n3502), .O(n3914) );
  FA1S U5006 ( .A(n3857), .B(n3856), .CI(n3855), .CO(n3926), .S(n3879) );
  XNR2HS U5007 ( .I1(n3931), .I2(n3930), .O(n3882) );
  FA1S U5008 ( .A(n3862), .B(n3861), .CI(n3860), .CO(n3945), .S(n3955) );
  FA1S U5009 ( .A(n3865), .B(n3864), .CI(n3863), .CO(n3846), .S(n3944) );
  FA1 U5010 ( .A(n3871), .B(n3870), .CI(n3869), .CO(n3845), .S(n3948) );
  FA1S U5011 ( .A(n3880), .B(n3879), .CI(n3878), .CO(n3931), .S(n3903) );
  MOAI1H U5012 ( .A1(n3901), .A2(n3881), .B1(n3903), .B2(n3902), .O(n3929) );
  XNR2HS U5013 ( .I1(n3882), .I2(n3929), .O(N6126) );
  INV1S U5014 ( .I(n61150), .O(n6084) );
  OAI12HS U5015 ( .B1(n6084), .B2(n6069), .A1(wait_conv_out_count[4]), .O(
        n3885) );
  NR2 U5016 ( .I1(N6291), .I2(wait_conv_out_count[1]), .O(n6094) );
  OAI12HS U5017 ( .B1(n6094), .B2(n3883), .A1(n5105), .O(n3884) );
  NR2 U5018 ( .I1(conv_temp[2]), .I2(product[2]), .O(n3886) );
  INV1S U5019 ( .I(image[7]), .O(n5609) );
  INV1S U5020 ( .I(image[6]), .O(n3900) );
  INV1S U5021 ( .I(image[5]), .O(n5606) );
  INV1S U5022 ( .I(image[4]), .O(n5605) );
  INV1S U5023 ( .I(image[3]), .O(n5604) );
  INV1S U5024 ( .I(image[2]), .O(n5603) );
  INV1S U5025 ( .I(n3902), .O(n3904) );
  XOR2HS U5026 ( .I1(n3904), .I2(n3903), .O(n3905) );
  XOR2HS U5027 ( .I1(n3901), .I2(n3905), .O(N6125) );
  XNR2HS U5028 ( .I1(n3907), .I2(n3906), .O(n3909) );
  XNR2HS U5029 ( .I1(n3909), .I2(n3908), .O(N6120) );
  NR2 U5030 ( .I1(n3509), .I2(n3495), .O(n3937) );
  NR2 U5031 ( .I1(n3910), .I2(n3495), .O(n3913) );
  NR2 U5032 ( .I1(n3509), .I2(n3500), .O(n3912) );
  NR2 U5033 ( .I1(n3510), .I2(n3495), .O(n3919) );
  NR2 U5034 ( .I1(n3509), .I2(n3502), .O(n3918) );
  NR2 U5035 ( .I1(n3910), .I2(n3500), .O(n3917) );
  FA1S U5036 ( .A(n3913), .B(n3912), .CI(n3911), .CO(n3936), .S(n3940) );
  FA1S U5037 ( .A(n3916), .B(n3915), .CI(n3914), .CO(n3925), .S(n3920) );
  FA1S U5038 ( .A(n3919), .B(n3918), .CI(n3917), .CO(n3911), .S(n3924) );
  FA1S U5039 ( .A(n3922), .B(n3921), .CI(n3920), .CO(n3923), .S(n3927) );
  FA1S U5040 ( .A(n3925), .B(n3924), .CI(n3923), .CO(n3939), .S(n3943) );
  FA1S U5041 ( .A(n3928), .B(n3927), .CI(n3926), .CO(n3942), .S(n3930) );
  INV1S U5042 ( .I(n3930), .O(n3934) );
  INV1S U5043 ( .I(n3931), .O(n3933) );
  OAI12H U5044 ( .B1(n3931), .B2(n3930), .A1(n3929), .O(n3932) );
  OAI12H U5045 ( .B1(n3934), .B2(n3933), .A1(n3932), .O(n3941) );
  FA1 U5046 ( .A(n3937), .B(n3936), .CI(n3935), .CO(N6130), .S(N6129) );
  FA1 U5047 ( .A(n3940), .B(n3939), .CI(n3938), .CO(n3935), .S(N6128) );
  FA1 U5048 ( .A(n3943), .B(n3942), .CI(n3941), .CO(n3938), .S(N6127) );
  FA1 U5049 ( .A(n3949), .B(n3948), .CI(n3947), .CO(n3974), .S(n3977) );
  FA1S U5050 ( .A(n3952), .B(n3951), .CI(n3950), .CO(n3976), .S(n3953) );
  FA1 U5051 ( .A(n3955), .B(n3954), .CI(n3953), .CO(n3979), .S(n3957) );
  ND2S U5052 ( .I1(n3980), .I2(n3979), .O(mult_x_231_n10) );
  NR2 U5053 ( .I1(n3979), .I2(n3980), .O(mult_x_231_n9) );
  FA1 U5054 ( .A(n3958), .B(n3957), .CI(n3956), .CO(mult_x_231_n11), .S(N6122)
         );
  FA1 U5055 ( .A(n3961), .B(n3960), .CI(n3959), .CO(n3956), .S(N6121) );
  FA1 U5056 ( .A(n3964), .B(n3963), .CI(n3962), .CO(n3908), .S(N6119) );
  FA1 U5057 ( .A(n3967), .B(n3966), .CI(n3965), .CO(n3962), .S(N6118) );
  FA1 U5058 ( .A(n3975), .B(n3974), .CI(n3973), .CO(n3902), .S(mult_x_231_n39)
         );
  NR2 U5059 ( .I1(n3515), .I2(n3494), .O(N6115) );
  INV1S U5060 ( .I(median_in[39]), .O(n5936) );
  INV1S U5061 ( .I(N1048), .O(n4040) );
  NR2 U5062 ( .I1(n4608), .I2(n4527), .O(n4018) );
  NR2 U5063 ( .I1(n5766), .I2(n3981), .O(n4046) );
  ND2S U5064 ( .I1(n4969), .I2(n6243), .O(n4098) );
  INV1S U5065 ( .I(n4098), .O(n4088) );
  ND2S U5066 ( .I1(n4046), .I2(n4088), .O(n3983) );
  ND3S U5067 ( .I1(n5725), .I2(n3537), .I3(n3992), .O(n4022) );
  AN2B1S U5068 ( .I1(n3984), .B1(n4606), .O(n3995) );
  NR2 U5069 ( .I1(n5010), .I2(n6245), .O(n4167) );
  INV1S U5070 ( .I(n4167), .O(n4055) );
  OAI12HS U5071 ( .B1(flip_flag), .B2(n5729), .A1(n3995), .O(n3985) );
  MOAI1S U5072 ( .A1(n4019), .A2(n4055), .B1(n5918), .B2(n3985), .O(n3990) );
  ND3S U5073 ( .I1(n4542), .I2(n4392), .I3(n5753), .O(n3988) );
  ND2S U5074 ( .I1(n3537), .I2(n3992), .O(n4021) );
  INV1S U5075 ( .I(n4021), .O(n3987) );
  INV1S U5076 ( .I(n4539), .O(n3986) );
  ND3S U5077 ( .I1(n3987), .I2(n5753), .I3(n3986), .O(n4026) );
  ND2S U5078 ( .I1(n3988), .I2(n4026), .O(n3989) );
  AOI22S U5079 ( .A1(n5755), .A2(n3990), .B1(n4025), .B2(n3989), .O(n3994) );
  NR2 U5080 ( .I1(n3992), .I2(n3993), .O(n5672) );
  NR2 U5081 ( .I1(state[1]), .I2(n3993), .O(n5670) );
  NR2 U5082 ( .I1(n5672), .I2(n5670), .O(n4358) );
  INV1S U5083 ( .I(n4358), .O(n4372) );
  NR2 U5084 ( .I1(n5744), .I2(n4372), .O(n4077) );
  INV1S U5085 ( .I(n6242), .O(n4599) );
  OAI12HS U5086 ( .B1(conv_sram_stop_flag_reg), .B2(n5669), .A1(n3537), .O(
        n5759) );
  INV3 U5087 ( .I(n5942), .O(n6064) );
  OAI112HS U5088 ( .C1(n3537), .C2(n4180), .A1(n4077), .B1(n6064), .O(n4035)
         );
  OAI112HS U5089 ( .C1(n4018), .C2(n4022), .A1(n3994), .B1(n4035), .O(n4371)
         );
  INV1S U5090 ( .I(n4371), .O(n5009) );
  INV1S U5091 ( .I(n5722), .O(n3997) );
  ND3S U5092 ( .I1(n4379), .I2(n5753), .I3(n4542), .O(n4032) );
  OAI22S U5093 ( .A1(n3997), .A2(n4032), .B1(n4034), .B2(n3996), .O(n4027) );
  NR2 U5094 ( .I1(image_size_temp[1]), .I2(cal_count[2]), .O(n3998) );
  NR2 U5095 ( .I1(n5746), .I2(n3998), .O(n4000) );
  AOI22S U5096 ( .A1(cal_count[2]), .A2(n3489), .B1(n3488), .B2(
        image_size_temp[1]), .O(n3999) );
  AN2S U5097 ( .I1(n5680), .I2(n4545), .O(n4037) );
  NR2 U5098 ( .I1(n4016), .I2(n4034), .O(n4010) );
  INV1S U5099 ( .I(cal_count_10[2]), .O(n5703) );
  INV1S U5100 ( .I(cal_count_10[1]), .O(n5708) );
  ND3S U5101 ( .I1(n5703), .I2(cal_count_10[3]), .I3(n5708), .O(n5696) );
  ND2S U5102 ( .I1(n4002), .I2(n5656), .O(n4008) );
  ND2S U5103 ( .I1(n4003), .I2(cal_count[1]), .O(n4006) );
  ND3S U5104 ( .I1(n4006), .I2(n4005), .I3(n4004), .O(n4007) );
  NR3 U5105 ( .I1(cal_count_10[0]), .I2(n5696), .I3(n4033), .O(n4013) );
  XOR2HS U5106 ( .I1(n4011), .I2(n5003), .O(n4999) );
  NR2 U5107 ( .I1(n4012), .I2(n4032), .O(n4028) );
  NR2 U5108 ( .I1(n4013), .I2(n4028), .O(n4015) );
  INV1S U5109 ( .I(cal_count_10[0]), .O(n5705) );
  NR2 U5110 ( .I1(n5708), .I2(n5705), .O(n5693) );
  ND2S U5111 ( .I1(n5693), .I2(n5703), .O(n5701) );
  OAI112HS U5112 ( .C1(n4016), .C2(n4034), .A1(n4015), .B1(n4014), .O(n4017)
         );
  XOR2HS U5113 ( .I1(n4017), .I2(n5003), .O(n4369) );
  INV1S U5114 ( .I(n4018), .O(n4023) );
  ND2S U5115 ( .I1(n5755), .I2(n4019), .O(n4020) );
  OAI12HS U5116 ( .B1(n4026), .B2(n4025), .A1(n4024), .O(n4036) );
  INV1S U5117 ( .I(n4036), .O(n4030) );
  NR2 U5118 ( .I1(n4028), .I2(n4027), .O(n4029) );
  ND2S U5119 ( .I1(n4030), .I2(n4029), .O(n4031) );
  ND3S U5120 ( .I1(n4034), .I2(n4033), .I3(n4032), .O(n4038) );
  OA13S U5121 ( .B1(n4038), .B2(n4037), .B3(n4036), .A1(n4035), .O(n5006) );
  MOAI1S U5122 ( .A1(n4040), .A2(n5009), .B1(n4039), .B2(n5006), .O(n2603) );
  INV1S U5123 ( .I(n4042), .O(n6131) );
  MOAI1S U5124 ( .A1(n4782), .A2(n6131), .B1(n4956), .B2(conv_temp[15]), .O(
        n2868) );
  INV1S U5125 ( .I(n4044), .O(n6132) );
  MOAI1S U5126 ( .A1(n4782), .A2(n6132), .B1(n4956), .B2(conv_temp[14]), .O(
        n2869) );
  INV1S U5127 ( .I(n4045), .O(n6241) );
  NR2 U5128 ( .I1(n4957), .I2(n6114), .O(n4947) );
  OAI112HS U5129 ( .C1(n6241), .C2(n4046), .A1(n4092), .B1(n4947), .O(n5558)
         );
  INV1S U5130 ( .I(n4180), .O(n5582) );
  NR2 U5131 ( .I1(state[0]), .I2(n4178), .O(n5677) );
  ND2S U5132 ( .I1(n5582), .I2(n5677), .O(n4076) );
  NR2 U5133 ( .I1(n5670), .I2(n5767), .O(n4179) );
  NR2 U5134 ( .I1(current_action_idx[1]), .I2(current_action_idx[2]), .O(n4169) );
  ND2S U5135 ( .I1(action_reg_2__2_), .I2(n4169), .O(n4048) );
  INV1S U5136 ( .I(current_action_idx[2]), .O(n4161) );
  NR2 U5137 ( .I1(current_action_idx[1]), .I2(n4161), .O(n4170) );
  INV1S U5138 ( .I(current_action_idx[1]), .O(n5662) );
  AOI22S U5139 ( .A1(n4170), .A2(action_reg_6__2_), .B1(n4171), .B2(
        action_reg_4__2_), .O(n4047) );
  ND3S U5140 ( .I1(n4048), .I2(n4047), .I3(current_action_idx[0]), .O(n4053)
         );
  ND2S U5141 ( .I1(action_reg_1__2_), .I2(n4169), .O(n4051) );
  AOI22S U5142 ( .A1(n4170), .A2(action_reg_5__2_), .B1(n4171), .B2(
        action_reg_3__2_), .O(n4050) );
  AOI13HS U5143 ( .B1(current_action_idx[2]), .B2(current_action_idx[1]), .B3(
        action_reg_7__2_), .A1(current_action_idx[0]), .O(n4049) );
  ND3S U5144 ( .I1(n4051), .I2(n4050), .I3(n4049), .O(n4052) );
  ND2S U5145 ( .I1(n4053), .I2(n4052), .O(n4363) );
  AO12S U5146 ( .B1(n4157), .B2(n4179), .A1(n4363), .O(n4054) );
  ND3S U5147 ( .I1(n4055), .I2(n4168), .I3(n4054), .O(n3405) );
  NR2 U5148 ( .I1(n4056), .I2(n3647), .O(n4166) );
  INV1S U5149 ( .I(image_size_reg[0]), .O(n61250) );
  ND2S U5150 ( .I1(image_size_reg[1]), .I2(n61250), .O(n4058) );
  ND2S U5151 ( .I1(SRAM_192X32_addr[4]), .I2(SRAM_192X32_addr[5]), .O(n4057)
         );
  NR2 U5152 ( .I1(n61250), .I2(image_size_reg[1]), .O(n4060) );
  NR2 U5153 ( .I1(SRAM_192X32_addr[4]), .I2(SRAM_192X32_addr[5]), .O(n4059) );
  MOAI1S U5154 ( .A1(n4058), .A2(n4057), .B1(n4060), .B2(n4059), .O(n4063) );
  OR3B2S U5155 ( .I1(n4060), .B1(n4059), .B2(n4058), .O(n4061) );
  NR3 U5156 ( .I1(n4061), .I2(SRAM_192X32_addr[2]), .I3(SRAM_192X32_addr[3]), 
        .O(n4062) );
  AO13S U5157 ( .B1(SRAM_192X32_addr[3]), .B2(SRAM_192X32_addr[2]), .B3(n4063), 
        .A1(n4062), .O(n4064) );
  AN3B2S U5158 ( .I1(SRAM_192X32_addr[7]), .B1(SRAM_192X32_addr[6]), .B2(n4065), .O(n4066) );
  MOAI1S U5159 ( .A1(state[0]), .A2(n3493), .B1(state[0]), .B2(n4066), .O(
        n4182) );
  ND3S U5160 ( .I1(n4069), .I2(n4068), .I3(n4067), .O(n5133) );
  AOI22S U5161 ( .A1(n4169), .A2(action_reg_2__0_), .B1(n4171), .B2(
        action_reg_4__0_), .O(n4075) );
  ND2S U5162 ( .I1(n4170), .I2(action_reg_6__0_), .O(n4074) );
  AOI22S U5163 ( .A1(n4170), .A2(action_reg_5__0_), .B1(n4171), .B2(
        action_reg_3__0_), .O(n4072) );
  ND2S U5164 ( .I1(n4169), .I2(action_reg_1__0_), .O(n4071) );
  ND3S U5165 ( .I1(current_action_idx[1]), .I2(current_action_idx[2]), .I3(
        action_reg_7__0_), .O(n4070) );
  AN4B1S U5166 ( .I1(n4072), .I2(n4071), .I3(n4070), .B1(current_action_idx[0]), .O(n4073) );
  AOI13HS U5167 ( .B1(current_action_idx[0]), .B2(n4075), .B3(n4074), .A1(
        n4073), .O(n4360) );
  ND2S U5168 ( .I1(n4077), .I2(n4076), .O(n4078) );
  MOAI1S U5169 ( .A1(n4182), .A2(n5133), .B1(n4360), .B2(n4078), .O(n4079) );
  NR2 U5170 ( .I1(n4166), .I2(n4079), .O(n4080) );
  INV1S U5171 ( .I(set_count[1]), .O(n5717) );
  INV1S U5172 ( .I(n5591), .O(n61230) );
  ND2S U5173 ( .I1(n61230), .I2(set_count[0]), .O(n5718) );
  NR2 U5174 ( .I1(n5717), .I2(n5718), .O(n5561) );
  ND2S U5175 ( .I1(set_count[2]), .I2(n5561), .O(n5557) );
  INV1S U5176 ( .I(SRAM_192_32_read_done), .O(n5668) );
  BUF6 U5177 ( .I(n4081), .O(n4743) );
  AOI22S U5178 ( .A1(n4193), .A2(SRAM_64X32_out_decode[0]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[24]), .O(n4085) );
  NR2 U5179 ( .I1(SRAM_192_32_read_done), .I2(n4082), .O(n4203) );
  NR2 U5180 ( .I1(n4542), .I2(n5668), .O(n4083) );
  BUF6 U5181 ( .I(n4083), .O(n4742) );
  AOI22S U5182 ( .A1(n3485), .A2(SRAM_192X32_out_decode[0]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[24]), .O(n4084) );
  ND2S U5183 ( .I1(n4085), .I2(n4084), .O(n4086) );
  MOAI1 U5184 ( .A1(n4748), .A2(n4086), .B1(n4748), .B2(n4086), .O(n5964) );
  ND3S U5185 ( .I1(n6243), .I2(n5725), .I3(n4623), .O(n5761) );
  NR2 U5186 ( .I1(n6064), .I2(n5761), .O(n4648) );
  MOAI1H U5187 ( .A1(n4623), .A2(n6064), .B1(n4648), .B2(n4191), .O(n4749) );
  AOI22S U5188 ( .A1(n4091), .A2(n4090), .B1(n4089), .B2(n5690), .O(n4383) );
  INV1S U5189 ( .I(n4092), .O(n4932) );
  OAI22S U5190 ( .A1(n4392), .A2(n4931), .B1(n4389), .B2(n4932), .O(n4093) );
  OAI22S U5191 ( .A1(n5751), .A2(n4512), .B1(n3486), .B2(n4512), .O(n4448) );
  AOI22S U5192 ( .A1(n5964), .A2(n4749), .B1(SRAM_out_buffer[24]), .B2(n4771), 
        .O(n4984) );
  NR2 U5193 ( .I1(n3486), .I2(n4381), .O(n4509) );
  ND3S U5194 ( .I1(n5656), .I2(cal_count[4]), .I3(cal_count[5]), .O(n4103) );
  NR3 U5195 ( .I1(n4945), .I2(n4094), .I3(n5749), .O(n5752) );
  NR2 U5196 ( .I1(n5751), .I2(n4096), .O(n4102) );
  INV1S U5197 ( .I(n5759), .O(n4386) );
  NR2 U5198 ( .I1(n5759), .I2(n3486), .O(n4375) );
  AOI13HS U5199 ( .B1(n5767), .B2(n4509), .B3(n5752), .A1(n4708), .O(n4688) );
  NR2 U5200 ( .I1(image_size_temp[1]), .I2(n6243), .O(n4380) );
  AOI22S U5201 ( .A1(n4388), .A2(n4932), .B1(n4380), .B2(n6309), .O(n4097) );
  NR2 U5202 ( .I1(n4097), .I2(n6064), .O(n4100) );
  AOI13HS U5203 ( .B1(n5753), .B2(n4098), .B3(n4386), .A1(n4100), .O(n4858) );
  INV1S U5204 ( .I(n4858), .O(n4099) );
  OAI12HS U5205 ( .B1(n4100), .B2(n4381), .A1(n4099), .O(n4432) );
  NR3 U5206 ( .I1(n3517), .I2(n5750), .I3(n4103), .O(n4104) );
  OAI22S U5207 ( .A1(n5752), .A2(n4393), .B1(n4394), .B2(n4104), .O(n4105) );
  AOI22S U5208 ( .A1(median_in[0]), .A2(n4981), .B1(median_in[8]), .B2(n6064), 
        .O(n4106) );
  NR2 U5209 ( .I1(n6245), .I2(n5756), .O(n4776) );
  INV1S U5210 ( .I(n4776), .O(n4894) );
  INV1S U5211 ( .I(n4894), .O(n4767) );
  INV1S U5212 ( .I(neg_flag), .O(n4746) );
  AOI22S U5213 ( .A1(n4743), .A2(SRAM_192X32_out_decode[28]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[28]), .O(n4108) );
  AOI22S U5214 ( .A1(n4193), .A2(SRAM_64X32_out_decode[4]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[4]), .O(n4107) );
  MOAI1 U5215 ( .A1(n5675), .A2(n4109), .B1(n5675), .B2(n4109), .O(n6044) );
  INV1S U5216 ( .I(n6044), .O(n5955) );
  AOI22S U5217 ( .A1(n5955), .A2(n4749), .B1(SRAM_out_buffer[28]), .B2(n4771), 
        .O(n5905) );
  AOI22S U5218 ( .A1(median_in[12]), .A2(n6064), .B1(median_in[4]), .B2(n4981), 
        .O(n4110) );
  INV1S U5219 ( .I(n4112), .O(n6134) );
  MOAI1S U5220 ( .A1(n4782), .A2(n6134), .B1(n4956), .B2(conv_temp[12]), .O(
        n2871) );
  INV1S U5221 ( .I(n4114), .O(n6133) );
  MOAI1S U5222 ( .A1(n4782), .A2(n6133), .B1(n4956), .B2(conv_temp[13]), .O(
        n2870) );
  BUF1 U5223 ( .I(n3487), .O(n6306) );
  BUF1 U5224 ( .I(n3487), .O(n6307) );
  FA1 U5225 ( .A(product[4]), .B(conv_temp[4]), .CI(n4115), .CO(n4121), .S(
        n4116) );
  INV1S U5226 ( .I(n4116), .O(n6142) );
  MOAI1S U5227 ( .A1(n4782), .A2(n6142), .B1(n4956), .B2(conv_temp[4]), .O(
        n2879) );
  INV1S U5228 ( .I(n4118), .O(n6144) );
  MOAI1S U5229 ( .A1(n4782), .A2(n6144), .B1(n4956), .B2(conv_temp[1]), .O(
        n2882) );
  XNR2HS U5230 ( .I1(product[2]), .I2(conv_temp[2]), .O(n4120) );
  MOAI1S U5231 ( .A1(n4782), .A2(n3504), .B1(n4956), .B2(conv_temp[2]), .O(
        n2881) );
  INV1S U5232 ( .I(n4122), .O(n6141) );
  MOAI1S U5233 ( .A1(n4782), .A2(n6141), .B1(n4956), .B2(conv_temp[5]), .O(
        n2878) );
  INV1S U5234 ( .I(n4124), .O(n6143) );
  MOAI1S U5235 ( .A1(n4782), .A2(n6143), .B1(n4956), .B2(conv_temp[3]), .O(
        n2880) );
  INV1S U5236 ( .I(n4125), .O(n61280) );
  MOAI1S U5237 ( .A1(n61280), .A2(n4782), .B1(n4956), .B2(conv_temp[0]), .O(
        n2883) );
  INV1S U5238 ( .I(n4127), .O(n6140) );
  MOAI1S U5239 ( .A1(n4782), .A2(n6140), .B1(n4956), .B2(conv_temp[6]), .O(
        n2877) );
  INV1S U5240 ( .I(SRAM_64X32_out_decode[10]), .O(n4128) );
  MOAI1S U5241 ( .A1(n6265), .A2(n4128), .B1(n6265), .B2(
        SRAM_64X32_data_out[10]), .O(n2642) );
  INV1S U5242 ( .I(SRAM_64X32_out_decode[20]), .O(n4129) );
  MOAI1S U5243 ( .A1(n6265), .A2(n4129), .B1(n6265), .B2(
        SRAM_64X32_data_out[20]), .O(n2685) );
  INV1S U5244 ( .I(SRAM_64X32_out_decode[11]), .O(n4130) );
  MOAI1S U5245 ( .A1(n6265), .A2(n4130), .B1(n6265), .B2(
        SRAM_64X32_data_out[11]), .O(n2651) );
  INV1S U5246 ( .I(SRAM_64X32_out_decode[2]), .O(n4131) );
  MOAI1S U5247 ( .A1(n6265), .A2(n4131), .B1(n6265), .B2(
        SRAM_64X32_data_out[2]), .O(n2684) );
  INV1S U5248 ( .I(SRAM_64X32_out_decode[17]), .O(n4132) );
  MOAI1S U5249 ( .A1(n6265), .A2(n4132), .B1(n6265), .B2(
        SRAM_64X32_data_out[17]), .O(n2681) );
  INV1S U5250 ( .I(SRAM_64X32_out_decode[19]), .O(n4133) );
  MOAI1S U5251 ( .A1(n6265), .A2(n4133), .B1(n6265), .B2(
        SRAM_64X32_data_out[19]), .O(n2683) );
  INV1S U5252 ( .I(SRAM_64X32_out_decode[16]), .O(n4134) );
  MOAI1S U5253 ( .A1(n6265), .A2(n4134), .B1(n6265), .B2(
        SRAM_64X32_data_out[16]), .O(n2680) );
  INV1S U5254 ( .I(SRAM_64X32_out_decode[1]), .O(n4135) );
  MOAI1S U5255 ( .A1(n6265), .A2(n4135), .B1(n6265), .B2(
        SRAM_64X32_data_out[1]), .O(n2633) );
  INV1S U5256 ( .I(SRAM_64X32_out_decode[12]), .O(n4136) );
  MOAI1S U5257 ( .A1(n6265), .A2(n4136), .B1(n6265), .B2(
        SRAM_64X32_data_out[12]), .O(n2660) );
  INV1S U5258 ( .I(SRAM_64X32_out_decode[15]), .O(n4137) );
  MOAI1S U5259 ( .A1(n6265), .A2(n4137), .B1(n6265), .B2(
        SRAM_64X32_data_out[15]), .O(n2679) );
  INV1S U5260 ( .I(SRAM_64X32_out_decode[18]), .O(n4138) );
  MOAI1S U5261 ( .A1(n6265), .A2(n4138), .B1(n6265), .B2(
        SRAM_64X32_data_out[18]), .O(n2682) );
  INV1S U5262 ( .I(SRAM_64X32_out_decode[13]), .O(n4139) );
  MOAI1S U5263 ( .A1(n6265), .A2(n4139), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_64X32_data_out[13]), .O(n2669) );
  INV1S U5264 ( .I(SRAM_64X32_out_decode[14]), .O(n4140) );
  MOAI1S U5265 ( .A1(n6265), .A2(n4140), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_64X32_data_out[14]), .O(n2678) );
  INV1S U5266 ( .I(SRAM_64X32_out_decode[7]), .O(n4141) );
  MOAI1S U5267 ( .A1(n6265), .A2(n4141), .B1(n6265), .B2(
        SRAM_64X32_data_out[7]), .O(n2701) );
  INV1S U5268 ( .I(SRAM_64X32_out_decode[6]), .O(n4142) );
  MOAI1S U5269 ( .A1(conv_sram_stop_flag_reg), .A2(n4142), .B1(
        conv_sram_stop_flag_reg), .B2(SRAM_64X32_data_out[6]), .O(n2700) );
  INV1S U5270 ( .I(SRAM_192X32_out_decode[17]), .O(n4143) );
  MOAI1S U5271 ( .A1(n6265), .A2(n4143), .B1(n6265), .B2(
        SRAM_192X32_data_out[17]), .O(n2721) );
  INV1S U5272 ( .I(SRAM_192X32_out_decode[16]), .O(n4144) );
  MOAI1S U5273 ( .A1(n6265), .A2(n4144), .B1(n6265), .B2(
        SRAM_192X32_data_out[16]), .O(n2720) );
  INV1S U5274 ( .I(SRAM_192X32_out_decode[22]), .O(n4145) );
  MOAI1S U5275 ( .A1(n6265), .A2(n4145), .B1(n6265), .B2(
        SRAM_192X32_data_out[22]), .O(n2727) );
  INV1S U5276 ( .I(SRAM_192X32_out_decode[21]), .O(n4146) );
  MOAI1S U5277 ( .A1(n6265), .A2(n4146), .B1(n6265), .B2(
        SRAM_192X32_data_out[21]), .O(n2726) );
  INV1S U5278 ( .I(SRAM_192X32_out_decode[25]), .O(n4147) );
  MOAI1S U5279 ( .A1(conv_sram_stop_flag_reg), .A2(n4147), .B1(n6265), .B2(
        SRAM_192X32_data_out[25]), .O(n2730) );
  INV1S U5280 ( .I(SRAM_192X32_out_decode[20]), .O(n4148) );
  MOAI1S U5281 ( .A1(conv_sram_stop_flag_reg), .A2(n4148), .B1(n6265), .B2(
        SRAM_192X32_data_out[20]), .O(n2725) );
  INV1S U5282 ( .I(SRAM_192X32_out_decode[19]), .O(n4149) );
  MOAI1S U5283 ( .A1(conv_sram_stop_flag_reg), .A2(n4149), .B1(n6265), .B2(
        SRAM_192X32_data_out[19]), .O(n2723) );
  INV1S U5284 ( .I(SRAM_192X32_out_decode[29]), .O(n4150) );
  MOAI1S U5285 ( .A1(conv_sram_stop_flag_reg), .A2(n4150), .B1(n6265), .B2(
        SRAM_192X32_data_out[29]), .O(n2734) );
  INV1S U5286 ( .I(SRAM_192X32_out_decode[28]), .O(n4151) );
  MOAI1S U5287 ( .A1(conv_sram_stop_flag_reg), .A2(n4151), .B1(n6265), .B2(
        SRAM_192X32_data_out[28]), .O(n2733) );
  INV1S U5288 ( .I(SRAM_192X32_out_decode[18]), .O(n4152) );
  MOAI1S U5289 ( .A1(n6265), .A2(n4152), .B1(n6265), .B2(
        SRAM_192X32_data_out[18]), .O(n2722) );
  INV1S U5290 ( .I(SRAM_192X32_out_decode[2]), .O(n4153) );
  MOAI1S U5291 ( .A1(n6265), .A2(n4153), .B1(n6265), .B2(
        SRAM_192X32_data_out[2]), .O(n2724) );
  INV1S U5292 ( .I(SRAM_192X32_out_decode[6]), .O(n4154) );
  MOAI1S U5293 ( .A1(conv_sram_stop_flag_reg), .A2(n4154), .B1(
        conv_sram_stop_flag_reg), .B2(SRAM_192X32_data_out[6]), .O(n2740) );
  FA1S U5294 ( .A(product[7]), .B(conv_temp[7]), .CI(n4155), .CO(n4162), .S(
        n4156) );
  INV1S U5295 ( .I(n4156), .O(n6139) );
  MOAI1S U5296 ( .A1(n4782), .A2(n6139), .B1(n4956), .B2(conv_temp[7]), .O(
        n2876) );
  INV1S U5297 ( .I(n4160), .O(n5665) );
  NR2 U5298 ( .I1(current_action_idx[0]), .I2(n5665), .O(n4158) );
  NR2 U5299 ( .I1(n61230), .I2(n4160), .O(n5661) );
  NR2 U5300 ( .I1(n4158), .I2(n5661), .O(n5663) );
  AO12S U5301 ( .B1(n4171), .B2(current_action_idx[0]), .A1(n4170), .O(n4159)
         );
  MOAI1S U5302 ( .A1(n5663), .A2(n4161), .B1(n4160), .B2(n4159), .O(n3230) );
  INV1S U5303 ( .I(n4163), .O(n6138) );
  MOAI1S U5304 ( .A1(n4782), .A2(n6138), .B1(n4956), .B2(conv_temp[8]), .O(
        n2875) );
  INV1S U5305 ( .I(n4165), .O(n6137) );
  MOAI1S U5306 ( .A1(n4782), .A2(n6137), .B1(n4956), .B2(conv_temp[9]), .O(
        n2874) );
  NR2 U5307 ( .I1(n4167), .I2(n4166), .O(n5013) );
  INV1S U5308 ( .I(n5712), .O(n4985) );
  AOI22S U5309 ( .A1(n4169), .A2(action_reg_2__1_), .B1(n4171), .B2(
        action_reg_4__1_), .O(n4177) );
  ND2S U5310 ( .I1(n4170), .I2(action_reg_6__1_), .O(n4176) );
  AOI22S U5311 ( .A1(n4170), .A2(action_reg_5__1_), .B1(n4169), .B2(
        action_reg_1__1_), .O(n4173) );
  ND2S U5312 ( .I1(action_reg_3__1_), .I2(n4171), .O(n4172) );
  OR3B2S U5313 ( .I1(current_action_idx[0]), .B1(n4173), .B2(n4172), .O(n4174)
         );
  AOI13HS U5314 ( .B1(current_action_idx[1]), .B2(current_action_idx[2]), .B3(
        action_reg_7__1_), .A1(n4174), .O(n4175) );
  AOI13HS U5315 ( .B1(current_action_idx[0]), .B2(n4177), .B3(n4176), .A1(
        n4175), .O(n4361) );
  ND2S U5316 ( .I1(n4179), .I2(n4178), .O(n4181) );
  AOI22S U5317 ( .A1(n4361), .A2(n4181), .B1(n5677), .B2(n4180), .O(n4184) );
  OR3B2S U5318 ( .I1(n5133), .B1(n4182), .B2(in_valid2), .O(n4183) );
  INV1S U5319 ( .I(n4186), .O(n6136) );
  MOAI1S U5320 ( .A1(n4782), .A2(n6136), .B1(n4956), .B2(conv_temp[10]), .O(
        n2873) );
  NR2 U5321 ( .I1(n4187), .I2(n5687), .O(n5655) );
  NR2 U5322 ( .I1(n5686), .I2(n5687), .O(n5659) );
  ND2S U5323 ( .I1(n3489), .I2(n5659), .O(n4188) );
  NR2 U5324 ( .I1(n5709), .I2(n4188), .O(n4189) );
  MOAI1S U5325 ( .A1(n4190), .A2(n5657), .B1(n4190), .B2(n4189), .O(n3234) );
  INV1S U5326 ( .I(n5766), .O(n4230) );
  OAI222S U5327 ( .A1(n4229), .A2(n4608), .B1(n4581), .B2(n4599), .C1(n4621), 
        .C2(n4230), .O(n4192) );
  AOI22S U5328 ( .A1(n4193), .A2(SRAM_64X32_out_decode[26]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[2]), .O(n4195) );
  AOI22S U5329 ( .A1(n3485), .A2(SRAM_192X32_out_decode[26]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[2]), .O(n4194) );
  ND2S U5330 ( .I1(n4195), .I2(n4194), .O(n4196) );
  MOAI1S U5331 ( .A1(n4748), .A2(n4196), .B1(n4748), .B2(n4196), .O(n5806) );
  INV2 U5332 ( .I(n5806), .O(n5867) );
  MOAI1S U5333 ( .A1(n5934), .A2(n5867), .B1(n5934), .B2(SRAM_out_buffer[66]), 
        .O(n3155) );
  AOI22S U5334 ( .A1(n4193), .A2(SRAM_64X32_out_decode[27]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[27]), .O(n4198) );
  AOI22S U5335 ( .A1(n4743), .A2(SRAM_192X32_out_decode[3]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[3]), .O(n4197) );
  MOAI1S U5336 ( .A1(n4746), .A2(n4199), .B1(n4746), .B2(n4199), .O(n5799) );
  INV1S U5337 ( .I(n5799), .O(n5870) );
  MOAI1S U5338 ( .A1(n5934), .A2(n5870), .B1(n5934), .B2(SRAM_out_buffer[67]), 
        .O(n3152) );
  AOI22S U5339 ( .A1(n3485), .A2(SRAM_192X32_out_decode[25]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[1]), .O(n4201) );
  AOI22S U5340 ( .A1(n4193), .A2(SRAM_64X32_out_decode[25]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[1]), .O(n4200) );
  ND2S U5341 ( .I1(n4201), .I2(n4200), .O(n4202) );
  MOAI1 U5342 ( .A1(n5675), .A2(n4202), .B1(n5675), .B2(n4202), .O(n5864) );
  MOAI1S U5343 ( .A1(n5934), .A2(n5864), .B1(n5934), .B2(SRAM_out_buffer[65]), 
        .O(n3158) );
  AOI22S U5344 ( .A1(n4193), .A2(SRAM_64X32_out_decode[21]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[13]), .O(n4205) );
  AOI22S U5345 ( .A1(n4203), .A2(SRAM_192X32_out_decode[21]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[13]), .O(n4204) );
  MOAI1 U5346 ( .A1(n5675), .A2(n4206), .B1(n5675), .B2(n4206), .O(n5875) );
  MOAI1S U5347 ( .A1(n5934), .A2(n5875), .B1(n5934), .B2(SRAM_out_buffer[77]), 
        .O(n3107) );
  INV1S U5348 ( .I(n4208), .O(n6135) );
  MOAI1S U5349 ( .A1(n4782), .A2(n6135), .B1(n4956), .B2(conv_temp[11]), .O(
        n2872) );
  INV1S U5350 ( .I(avg_temp[4]), .O(n6285) );
  NR2 U5351 ( .I1(avg_temp[8]), .I2(n4210), .O(n6198) );
  INV1S U5352 ( .I(n6198), .O(n4211) );
  ND2S U5353 ( .I1(n4211), .I2(n4212), .O(n6199) );
  MOAI1S U5354 ( .A1(avg_temp[7]), .A2(n6198), .B1(avg_temp[7]), .B2(n6199), 
        .O(n4213) );
  INV1S U5355 ( .I(avg_temp[7]), .O(n6273) );
  AOI22S U5356 ( .A1(n6273), .A2(n4212), .B1(avg_temp[7]), .B2(n4211), .O(
        n4226) );
  INV1S U5357 ( .I(avg_temp[6]), .O(n6277) );
  NR2 U5358 ( .I1(n6277), .I2(n4213), .O(n4227) );
  MOAI1S U5359 ( .A1(avg_temp[6]), .A2(n4226), .B1(avg_temp[6]), .B2(n4226), 
        .O(n4214) );
  NR2 U5360 ( .I1(n4227), .I2(n4214), .O(n4218) );
  OR2B1S U5361 ( .I1(n4216), .B1(n4215), .O(n6202) );
  OAI12HS U5362 ( .B1(avg_temp[5]), .B2(n4216), .A1(n4217), .O(n4221) );
  NR2 U5363 ( .I1(n6285), .I2(n4221), .O(n4219) );
  INV1S U5364 ( .I(avg_temp[5]), .O(n6281) );
  MOAI1S U5365 ( .A1(n4218), .A2(n4217), .B1(n4218), .B2(n6281), .O(n4224) );
  NR2 U5366 ( .I1(n4219), .I2(n4224), .O(n4220) );
  MOAI1S U5367 ( .A1(n6219), .A2(n4220), .B1(n6219), .B2(gray_avg_reg[28]), 
        .O(n2772) );
  NR2 U5368 ( .I1(n4220), .I2(n6285), .O(n4222) );
  MOAI1S U5369 ( .A1(n4221), .A2(avg_temp[4]), .B1(n4221), .B2(n4222), .O(
        n4869) );
  INV1S U5370 ( .I(n4222), .O(n4223) );
  OAI22S U5371 ( .A1(avg_temp[3]), .A2(n4869), .B1(n4871), .B2(n4869), .O(
        n4225) );
  MOAI1S U5372 ( .A1(n6219), .A2(n4225), .B1(n6219), .B2(gray_avg_reg[27]), 
        .O(n2771) );
  NR2 U5373 ( .I1(n4227), .I2(n4226), .O(n4228) );
  MOAI1S U5374 ( .A1(n6219), .A2(n4228), .B1(n6219), .B2(gray_avg_reg[30]), 
        .O(n2774) );
  INV1S U5375 ( .I(n4229), .O(n5763) );
  MOAI1S U5376 ( .A1(n4230), .A2(n4608), .B1(n5758), .B2(n5763), .O(n4231) );
  NR2 U5377 ( .I1(n4623), .I2(n6064), .O(n4647) );
  AOI22S U5378 ( .A1(n4743), .A2(SRAM_192X32_out_decode[11]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[11]), .O(n4233) );
  AOI22S U5379 ( .A1(n4193), .A2(SRAM_64X32_out_decode[19]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[19]), .O(n4232) );
  MOAI1 U5380 ( .A1(n5675), .A2(n4234), .B1(n5675), .B2(n4234), .O(n5869) );
  MOAI1S U5381 ( .A1(n5933), .A2(n5869), .B1(n5933), .B2(SRAM_out_buffer[43]), 
        .O(n3120) );
  MOAI1S U5382 ( .A1(n5933), .A2(n5875), .B1(n5933), .B2(SRAM_out_buffer[45]), 
        .O(n3108) );
  AOI22S U5383 ( .A1(n4193), .A2(SRAM_64X32_out_decode[18]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[10]), .O(n4236) );
  AOI22S U5384 ( .A1(n3485), .A2(SRAM_192X32_out_decode[18]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[10]), .O(n4235) );
  MOAI1 U5385 ( .A1(n5675), .A2(n4237), .B1(n5675), .B2(n4237), .O(n5866) );
  MOAI1S U5386 ( .A1(n5933), .A2(n5866), .B1(n5933), .B2(SRAM_out_buffer[42]), 
        .O(n3126) );
  AOI22S U5387 ( .A1(n3485), .A2(SRAM_192X32_out_decode[22]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[14]), .O(n4239) );
  AOI22S U5388 ( .A1(n4193), .A2(SRAM_64X32_out_decode[22]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[14]), .O(n4238) );
  MOAI1 U5389 ( .A1(n5675), .A2(n4240), .B1(n5675), .B2(n4240), .O(n5878) );
  MOAI1S U5390 ( .A1(n5933), .A2(n5878), .B1(n5933), .B2(SRAM_out_buffer[46]), 
        .O(n3102) );
  AOI22S U5391 ( .A1(n4743), .A2(SRAM_192X32_out_decode[8]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[8]), .O(n4242) );
  AOI22S U5392 ( .A1(n4193), .A2(SRAM_64X32_out_decode[16]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[16]), .O(n4241) );
  ND2S U5393 ( .I1(n4242), .I2(n4241), .O(n4243) );
  MOAI1S U5394 ( .A1(n4748), .A2(n4243), .B1(n4748), .B2(n4243), .O(n5805) );
  MOAI1S U5395 ( .A1(n5933), .A2(n5860), .B1(n5933), .B2(SRAM_out_buffer[40]), 
        .O(n3138) );
  AOI22S U5396 ( .A1(n4193), .A2(SRAM_64X32_out_decode[29]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[5]), .O(n4245) );
  AOI22S U5397 ( .A1(n3485), .A2(SRAM_192X32_out_decode[29]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[5]), .O(n4244) );
  MOAI1S U5398 ( .A1(n4746), .A2(n4246), .B1(n4748), .B2(n4246), .O(n5791) );
  INV1S U5399 ( .I(n5791), .O(n5876) );
  MOAI1S U5400 ( .A1(n5933), .A2(n5876), .B1(n5933), .B2(SRAM_out_buffer[37]), 
        .O(n3147) );
  AOI22S U5401 ( .A1(SRAM_192X32_out_decode[9]), .A2(n4743), .B1(
        SRAM_64X32_out_decode[9]), .B2(n4742), .O(n4248) );
  AOI22S U5402 ( .A1(SRAM_64X32_out_decode[17]), .A2(n4193), .B1(
        SRAM_192X32_out_decode[17]), .B2(n3485), .O(n4247) );
  MOAI1S U5403 ( .A1(n4748), .A2(n4249), .B1(n4748), .B2(n4249), .O(n5804) );
  INV2 U5404 ( .I(n5804), .O(n5863) );
  MOAI1S U5405 ( .A1(n5933), .A2(n5863), .B1(n5933), .B2(SRAM_out_buffer[41]), 
        .O(n3132) );
  AOI22S U5406 ( .A1(n3485), .A2(SRAM_192X32_out_decode[30]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[6]), .O(n4251) );
  AOI22S U5407 ( .A1(n4193), .A2(SRAM_64X32_out_decode[30]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[6]), .O(n4250) );
  MOAI1S U5408 ( .A1(n4748), .A2(n4252), .B1(n4748), .B2(n4252), .O(n5813) );
  INV1S U5409 ( .I(n5813), .O(n5881) );
  MOAI1S U5410 ( .A1(n5933), .A2(n5881), .B1(n5933), .B2(SRAM_out_buffer[38]), 
        .O(n3144) );
  AOI22S U5411 ( .A1(n4193), .A2(SRAM_64X32_out_decode[15]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[23]), .O(n4254) );
  AOI22S U5412 ( .A1(n3485), .A2(SRAM_192X32_out_decode[15]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[23]), .O(n4253) );
  MOAI1S U5413 ( .A1(n4748), .A2(n4255), .B1(n4748), .B2(n4255), .O(n5969) );
  INV1S U5414 ( .I(n5969), .O(n6029) );
  MOAI1S U5415 ( .A1(n5933), .A2(n6029), .B1(n5933), .B2(SRAM_out_buffer[55]), 
        .O(n3016) );
  MOAI1S U5416 ( .A1(n5933), .A2(n5864), .B1(n5933), .B2(SRAM_out_buffer[33]), 
        .O(n3159) );
  AOI22S U5417 ( .A1(n4193), .A2(SRAM_64X32_out_decode[23]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[15]), .O(n4257) );
  AOI22S U5418 ( .A1(n3485), .A2(SRAM_192X32_out_decode[23]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[15]), .O(n4256) );
  MOAI1 U5419 ( .A1(n5675), .A2(n4258), .B1(n5675), .B2(n4258), .O(n5857) );
  MOAI1S U5420 ( .A1(n5933), .A2(n5857), .B1(n5933), .B2(SRAM_out_buffer[47]), 
        .O(n3096) );
  AOI22S U5421 ( .A1(n4743), .A2(SRAM_192X32_out_decode[18]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[18]), .O(n4260) );
  AOI22S U5422 ( .A1(n4193), .A2(SRAM_64X32_out_decode[10]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[10]), .O(n4259) );
  MOAI1 U5423 ( .A1(n5675), .A2(n4261), .B1(n5675), .B2(n4261), .O(n6037) );
  MOAI1S U5424 ( .A1(n5933), .A2(n6037), .B1(n5933), .B2(SRAM_out_buffer[50]), 
        .O(n3046) );
  INV1S U5425 ( .I(median_in[15]), .O(n6067) );
  INV1S U5426 ( .I(median_in[7]), .O(n5276) );
  NR2 U5427 ( .I1(n5276), .I2(median_in[23]), .O(n5255) );
  NR2 U5428 ( .I1(median_in[7]), .I2(n6067), .O(n5223) );
  INV1S U5429 ( .I(median_in[23]), .O(n5275) );
  NR2 U5430 ( .I1(median_in[7]), .I2(n5275), .O(n5243) );
  NR2 U5431 ( .I1(n5223), .I2(n5243), .O(n4785) );
  INV1S U5432 ( .I(median_in[14]), .O(n5270) );
  AOI22S U5433 ( .A1(median_in[22]), .A2(n5270), .B1(median_in[23]), .B2(n6067), .O(n5232) );
  INV1S U5434 ( .I(median_in[9]), .O(n5263) );
  AOI22S U5435 ( .A1(median_in[17]), .A2(n5263), .B1(median_in[18]), .B2(n5265), .O(n5227) );
  INV1S U5436 ( .I(median_in[16]), .O(n5260) );
  MOAI1S U5437 ( .A1(median_in[17]), .A2(n5263), .B1(n5260), .B2(median_in[8]), 
        .O(n4262) );
  OAI22S U5438 ( .A1(n5227), .A2(n5226), .B1(n4262), .B2(n5226), .O(n4266) );
  INV1S U5439 ( .I(median_in[11]), .O(n5267) );
  INV1S U5440 ( .I(median_in[12]), .O(n5906) );
  AOI22S U5441 ( .A1(median_in[19]), .A2(n5267), .B1(median_in[20]), .B2(n5906), .O(n4263) );
  INV1S U5442 ( .I(median_in[13]), .O(n5922) );
  MOAI1S U5443 ( .A1(median_in[22]), .A2(n5270), .B1(n5919), .B2(median_in[13]), .O(n4264) );
  AOI13HS U5444 ( .B1(median_in[12]), .B2(n4265), .B3(n5909), .A1(n4264), .O(
        n5228) );
  OAI12HS U5445 ( .B1(n4266), .B2(n5229), .A1(n5228), .O(n4267) );
  MOAI1S U5446 ( .A1(n5259), .A2(median_in[14]), .B1(n5259), .B2(n5271), .O(
        n4276) );
  MOAI1S U5447 ( .A1(n5259), .A2(median_in[13]), .B1(n5259), .B2(n5919), .O(
        n5278) );
  MOAI1S U5448 ( .A1(n5259), .A2(median_in[12]), .B1(n5259), .B2(n5909), .O(
        n4277) );
  MOAI1S U5449 ( .A1(n5259), .A2(median_in[11]), .B1(n5259), .B2(n5268), .O(
        n4278) );
  INV1S U5450 ( .I(median_in[18]), .O(n5266) );
  MOAI1S U5451 ( .A1(n5259), .A2(median_in[10]), .B1(n5259), .B2(n5266), .O(
        n4275) );
  FA1S U5452 ( .A(median_in[1]), .B(n5277), .CI(n4274), .CO(n4268) );
  FA1S U5453 ( .A(n4275), .B(median_in[2]), .CI(n4268), .CO(n4269) );
  FA1S U5454 ( .A(median_in[3]), .B(n4278), .CI(n4269), .CO(n4270) );
  MOAI1S U5455 ( .A1(n5279), .A2(n4274), .B1(n5279), .B2(median_in[1]), .O(
        find_median_inst_max3[1]) );
  MOAI1S U5456 ( .A1(n5279), .A2(n4275), .B1(n5279), .B2(median_in[2]), .O(
        find_median_inst_max3[2]) );
  MOAI1S U5457 ( .A1(n5279), .A2(n4276), .B1(n5279), .B2(median_in[6]), .O(
        find_median_inst_max3[6]) );
  MOAI1S U5458 ( .A1(n5279), .A2(n4277), .B1(n5279), .B2(median_in[4]), .O(
        find_median_inst_max3[4]) );
  MOAI1S U5459 ( .A1(n5279), .A2(n4278), .B1(n5279), .B2(median_in[3]), .O(
        find_median_inst_max3[3]) );
  NR2 U5460 ( .I1(median_in[39]), .I2(median_in[47]), .O(n4292) );
  INV1S U5461 ( .I(median_in[34]), .O(n5178) );
  AOI22S U5462 ( .A1(median_in[43]), .A2(n5890), .B1(median_in[42]), .B2(n5178), .O(n5142) );
  OAI22S U5463 ( .A1(median_in[41]), .A2(median_in[40]), .B1(n5177), .B2(
        median_in[40]), .O(n5144) );
  INV1S U5464 ( .I(median_in[43]), .O(n5186) );
  AOI22S U5465 ( .A1(n5142), .A2(n4279), .B1(median_in[35]), .B2(n5186), .O(
        n4284) );
  INV1S U5466 ( .I(median_in[46]), .O(n5183) );
  NR2 U5467 ( .I1(median_in[38]), .I2(n5183), .O(n4283) );
  INV1S U5468 ( .I(median_in[37]), .O(n5910) );
  NR2 U5469 ( .I1(median_in[45]), .I2(n5910), .O(n4281) );
  INV1S U5470 ( .I(median_in[44]), .O(n5185) );
  AOI13HS U5471 ( .B1(median_in[36]), .B2(n5185), .B3(n4282), .A1(n4281), .O(
        n5148) );
  OAI22S U5472 ( .A1(n4284), .A2(n5145), .B1(n4283), .B2(n5148), .O(n4285) );
  INV1S U5473 ( .I(median_in[38]), .O(n5923) );
  MOAI1S U5474 ( .A1(median_in[46]), .A2(n5923), .B1(n5205), .B2(median_in[39]), .O(n5149) );
  OAI22H U5475 ( .A1(n4285), .A2(n5149), .B1(n5205), .B2(median_in[39]), .O(
        n5187) );
  MOAI1S U5476 ( .A1(n5208), .A2(median_in[46]), .B1(n5208), .B2(n5923), .O(
        n4294) );
  MOAI1S U5477 ( .A1(n5208), .A2(median_in[45]), .B1(n5208), .B2(n5910), .O(
        n5210) );
  INV1S U5478 ( .I(median_in[36]), .O(n5899) );
  MOAI1S U5479 ( .A1(n5208), .A2(median_in[44]), .B1(n5208), .B2(n5899), .O(
        n4295) );
  MOAI1S U5480 ( .A1(n5208), .A2(median_in[43]), .B1(n5208), .B2(n5890), .O(
        n4297) );
  MOAI1S U5481 ( .A1(n5208), .A2(median_in[42]), .B1(n5208), .B2(n5178), .O(
        n4293) );
  FA1S U5482 ( .A(median_in[25]), .B(median_in[24]), .CI(n4296), .CO(n4286) );
  FA1S U5483 ( .A(median_in[26]), .B(n4293), .CI(n4286), .CO(n4287) );
  FA1S U5484 ( .A(n4297), .B(median_in[27]), .CI(n4287), .CO(n4288) );
  FA1S U5485 ( .A(median_in[28]), .B(n4295), .CI(n4288), .CO(n4289) );
  MOAI1S U5486 ( .A1(n5211), .A2(n4293), .B1(n5211), .B2(median_in[26]), .O(
        find_median_inst_max2[2]) );
  MOAI1S U5487 ( .A1(n5211), .A2(n4294), .B1(n5211), .B2(median_in[30]), .O(
        find_median_inst_max2[6]) );
  MOAI1S U5488 ( .A1(n5211), .A2(n4295), .B1(n5211), .B2(median_in[28]), .O(
        find_median_inst_max2[4]) );
  MOAI1S U5489 ( .A1(n5211), .A2(n4296), .B1(n5211), .B2(median_in[25]), .O(
        find_median_inst_max2[1]) );
  MOAI1S U5490 ( .A1(n5211), .A2(n4297), .B1(n5211), .B2(median_in[27]), .O(
        find_median_inst_max2[3]) );
  MOAI1S U5491 ( .A1(n5233), .A2(median_in[14]), .B1(n5233), .B2(n5271), .O(
        n4306) );
  MOAI1S U5492 ( .A1(n5233), .A2(median_in[13]), .B1(n5233), .B2(n5919), .O(
        n4311) );
  MOAI1S U5493 ( .A1(n5259), .A2(median_in[20]), .B1(n5259), .B2(n5906), .O(
        n4308) );
  MOAI1S U5494 ( .A1(n5233), .A2(median_in[11]), .B1(n5233), .B2(n5268), .O(
        n4310) );
  MOAI1S U5495 ( .A1(n5233), .A2(median_in[10]), .B1(n5233), .B2(n5266), .O(
        n4309) );
  FA1S U5496 ( .A(median_in[1]), .B(median_in[0]), .CI(n4307), .CO(n4298) );
  FA1S U5497 ( .A(n4309), .B(median_in[2]), .CI(n4298), .CO(n4299) );
  FA1S U5498 ( .A(median_in[3]), .B(n4310), .CI(n4299), .CO(n4300) );
  FA1S U5499 ( .A(n4308), .B(median_in[4]), .CI(n4300), .CO(n4301) );
  NR2 U5500 ( .I1(n5276), .I2(median_in[15]), .O(n5221) );
  MOAI1S U5501 ( .A1(n5233), .A2(median_in[8]), .B1(n5233), .B2(n5260), .O(
        n4305) );
  MOAI1S U5502 ( .A1(n4312), .A2(n4305), .B1(n4312), .B2(median_in[0]), .O(
        find_median_inst_min3[0]) );
  MOAI1S U5503 ( .A1(n4312), .A2(n4306), .B1(n4312), .B2(median_in[6]), .O(
        find_median_inst_min3[6]) );
  MOAI1S U5504 ( .A1(n4312), .A2(n4307), .B1(n4312), .B2(median_in[1]), .O(
        find_median_inst_min3[1]) );
  MOAI1S U5505 ( .A1(n4312), .A2(n4308), .B1(n4312), .B2(median_in[4]), .O(
        find_median_inst_min3[4]) );
  MOAI1S U5506 ( .A1(n4312), .A2(n4309), .B1(n4312), .B2(median_in[2]), .O(
        find_median_inst_min3[2]) );
  MOAI1S U5507 ( .A1(n4312), .A2(n4310), .B1(n4312), .B2(median_in[3]), .O(
        find_median_inst_min3[3]) );
  MOAI1S U5508 ( .A1(n4312), .A2(n4311), .B1(n4312), .B2(median_in[5]), .O(
        find_median_inst_min3[5]) );
  INV1S U5509 ( .I(median_in[71]), .O(n5945) );
  INV1S U5510 ( .I(median_in[55]), .O(n5940) );
  INV1S U5511 ( .I(n5542), .O(n5499) );
  INV1S U5512 ( .I(median_in[63]), .O(n5944) );
  NR2 U5513 ( .I1(median_in[55]), .I2(n5944), .O(n5504) );
  NR2 U5514 ( .I1(n5499), .I2(n5504), .O(n4784) );
  INV1S U5515 ( .I(median_in[62]), .O(n5928) );
  MOAI1S U5516 ( .A1(median_in[70]), .A2(n5928), .B1(n5945), .B2(median_in[63]), .O(n5496) );
  NR2 U5517 ( .I1(median_in[62]), .I2(n5927), .O(n4319) );
  NR2 U5518 ( .I1(median_in[69]), .I2(n5914), .O(n4314) );
  AOI13HS U5519 ( .B1(median_in[60]), .B2(n5532), .B3(n4315), .A1(n4314), .O(
        n5495) );
  INV1S U5520 ( .I(median_in[56]), .O(n5524) );
  MOAI1S U5521 ( .A1(median_in[64]), .A2(n5524), .B1(n5534), .B2(median_in[57]), .O(n4313) );
  ND2S U5522 ( .I1(median_in[65]), .I2(n5525), .O(n5485) );
  INV1S U5523 ( .I(median_in[58]), .O(n5527) );
  ND2S U5524 ( .I1(median_in[66]), .I2(n5527), .O(n5491) );
  INV1S U5525 ( .I(median_in[66]), .O(n5533) );
  AOI13HS U5526 ( .B1(n4317), .B2(n5494), .B3(n5487), .A1(n5492), .O(n4318) );
  INV1S U5527 ( .I(median_in[59]), .O(n5895) );
  MOAI1S U5528 ( .A1(n5546), .A2(median_in[70]), .B1(n5546), .B2(n5928), .O(
        n5555) );
  INV1S U5529 ( .I(median_in[69]), .O(n5913) );
  MOAI1S U5530 ( .A1(n5520), .A2(median_in[61]), .B1(n5520), .B2(n5913), .O(
        n4328) );
  INV1S U5531 ( .I(median_in[60]), .O(n5902) );
  MOAI1S U5532 ( .A1(n5546), .A2(median_in[68]), .B1(n5546), .B2(n5902), .O(
        n4330) );
  MOAI1S U5533 ( .A1(n5546), .A2(median_in[67]), .B1(n5546), .B2(n5895), .O(
        n4329) );
  MOAI1S U5534 ( .A1(n5546), .A2(median_in[66]), .B1(n5546), .B2(n5527), .O(
        n4327) );
  FA1S U5535 ( .A(median_in[49]), .B(median_in[48]), .CI(n4332), .CO(n4321) );
  FA1S U5536 ( .A(median_in[50]), .B(n4327), .CI(n4321), .CO(n4322) );
  FA1S U5537 ( .A(n4329), .B(median_in[51]), .CI(n4322), .CO(n4323) );
  MOAI1S U5538 ( .A1(n5556), .A2(n4327), .B1(n5556), .B2(median_in[50]), .O(
        find_median_inst_max1[2]) );
  MOAI1S U5539 ( .A1(n5556), .A2(n4328), .B1(n5556), .B2(median_in[53]), .O(
        find_median_inst_max1[5]) );
  MOAI1S U5540 ( .A1(n5556), .A2(n4329), .B1(n5556), .B2(median_in[51]), .O(
        find_median_inst_max1[3]) );
  MOAI1S U5541 ( .A1(n5556), .A2(n4330), .B1(n5556), .B2(median_in[52]), .O(
        find_median_inst_max1[4]) );
  INV1S U5542 ( .I(median_in[64]), .O(n5545) );
  MOAI1S U5543 ( .A1(n5520), .A2(median_in[56]), .B1(n5520), .B2(n5545), .O(
        n4331) );
  MOAI1S U5544 ( .A1(n5556), .A2(n4331), .B1(n5556), .B2(median_in[48]), .O(
        find_median_inst_max1[0]) );
  MOAI1S U5545 ( .A1(n5556), .A2(n4332), .B1(n5556), .B2(median_in[49]), .O(
        find_median_inst_max1[1]) );
  NR2 U5546 ( .I1(find_median_inst_min1_reg[7]), .I2(
        find_median_inst_min2_reg[7]), .O(n4355) );
  INV1S U5547 ( .I(find_median_inst_min2_reg[7]), .O(n4345) );
  INV1S U5548 ( .I(find_median_inst_min2_reg[6]), .O(n4343) );
  INV1S U5549 ( .I(find_median_inst_min2_reg[5]), .O(n4341) );
  INV1S U5550 ( .I(find_median_inst_min2_reg[4]), .O(n4339) );
  INV1S U5551 ( .I(find_median_inst_min2_reg[3]), .O(n4337) );
  INV1S U5552 ( .I(find_median_inst_min2_reg[2]), .O(n4335) );
  INV1S U5553 ( .I(find_median_inst_min2_reg[1]), .O(n4333) );
  OAI22S U5554 ( .A1(n4347), .A2(find_median_inst_min1_reg[6]), .B1(n4346), 
        .B2(find_median_inst_min2_reg[6]), .O(n5396) );
  OAI22S U5555 ( .A1(n4347), .A2(find_median_inst_min1_reg[5]), .B1(n4346), 
        .B2(find_median_inst_min2_reg[5]), .O(n5395) );
  OAI22S U5556 ( .A1(n4347), .A2(find_median_inst_min1_reg[4]), .B1(n4346), 
        .B2(find_median_inst_min2_reg[4]), .O(n5394) );
  OAI22S U5557 ( .A1(n4347), .A2(find_median_inst_min1_reg[3]), .B1(n4346), 
        .B2(find_median_inst_min2_reg[3]), .O(n5393) );
  OAI22S U5558 ( .A1(n4347), .A2(find_median_inst_min1_reg[2]), .B1(n4346), 
        .B2(find_median_inst_min2_reg[2]), .O(n5392) );
  OAI22S U5559 ( .A1(n4346), .A2(find_median_inst_min2_reg[0]), .B1(n4347), 
        .B2(find_median_inst_min1_reg[0]), .O(n4354) );
  OAI22S U5560 ( .A1(n4347), .A2(find_median_inst_min1_reg[1]), .B1(n4346), 
        .B2(find_median_inst_min2_reg[1]), .O(n5391) );
  MOAI1S U5561 ( .A1(n5397), .A2(n4354), .B1(n5397), .B2(
        find_median_inst_min3_reg[0]), .O(find_median_inst_min_max[0]) );
  OR2B1S U5562 ( .I1(find_median_inst_min3_reg[7]), .B1(n4355), .O(
        find_median_inst_min_max[7]) );
  ND2S U5563 ( .I1(n4357), .I2(n5006), .O(n4367) );
  ND2S U5564 ( .I1(n4371), .I2(N1043), .O(n4366) );
  INV1S U5565 ( .I(n4547), .O(n4598) );
  ND2S U5566 ( .I1(state[0]), .I2(n5670), .O(n4359) );
  MOAI1S U5567 ( .A1(flip_flag), .A2(n4359), .B1(flip_flag), .B2(n4359), .O(
        n5590) );
  ND3S U5568 ( .I1(n4361), .I2(n5590), .I3(n4360), .O(n4362) );
  NR2 U5569 ( .I1(n4363), .I2(n4362), .O(n5068) );
  ND3S U5570 ( .I1(n5068), .I2(n5766), .I3(n5682), .O(n4364) );
  NR2 U5571 ( .I1(n4598), .I2(n4364), .O(n5125) );
  INV1S U5572 ( .I(n5125), .O(n4365) );
  FA1S U5573 ( .A(N1044), .B(n4369), .CI(n4368), .CO(n4998), .S(n4370) );
  ND2S U5574 ( .I1(n4370), .I2(n5006), .O(n4374) );
  ND2S U5575 ( .I1(n4371), .I2(N1044), .O(n4373) );
  ND3S U5576 ( .I1(n4372), .I2(n5068), .I3(n5755), .O(n5109) );
  OAI112HS U5577 ( .C1(image_size_temp[1]), .C2(n4376), .A1(n4386), .B1(n6309), 
        .O(n4377) );
  OAI22S U5578 ( .A1(n4379), .A2(n4391), .B1(n4378), .B2(n4377), .O(n4466) );
  ND2S U5579 ( .I1(SRAM_out_buffer[65]), .I2(n4466), .O(n4397) );
  OAI12HS U5580 ( .B1(n4381), .B2(n6309), .A1(n4380), .O(n4382) );
  AO13S U5581 ( .B1(n4383), .B2(n4382), .B3(n4387), .A1(n5918), .O(n4384) );
  ND2 U5582 ( .I1(n5942), .I2(n4384), .O(n4385) );
  ND3S U5583 ( .I1(n4388), .I2(n4387), .I3(n4386), .O(n4390) );
  OAI22S U5584 ( .A1(n4392), .A2(n4391), .B1(n4390), .B2(n4389), .O(n5770) );
  AOI22S U5585 ( .A1(window_1__4__1_), .A2(n4385), .B1(SRAM_out_buffer[33]), 
        .B2(n4416), .O(n4396) );
  INV1S U5586 ( .I(n4510), .O(n4709) );
  AOI22S U5587 ( .A1(SRAM_out_buffer[41]), .A2(n4709), .B1(SRAM_out_buffer[73]), .B2(n4708), .O(n4395) );
  ND2S U5588 ( .I1(SRAM_out_buffer[64]), .I2(n4466), .O(n4400) );
  AOI22S U5589 ( .A1(window_1__4__0_), .A2(n4385), .B1(SRAM_out_buffer[32]), 
        .B2(n4416), .O(n4399) );
  AOI22S U5590 ( .A1(SRAM_out_buffer[40]), .A2(n4709), .B1(SRAM_out_buffer[72]), .B2(n4708), .O(n4398) );
  ND2S U5591 ( .I1(SRAM_out_buffer[66]), .I2(n4466), .O(n4403) );
  AOI22S U5592 ( .A1(window_1__4__2_), .A2(n4385), .B1(SRAM_out_buffer[34]), 
        .B2(n4416), .O(n4402) );
  AOI22S U5593 ( .A1(SRAM_out_buffer[42]), .A2(n4709), .B1(SRAM_out_buffer[74]), .B2(n4708), .O(n4401) );
  ND2S U5594 ( .I1(SRAM_out_buffer[69]), .I2(n4466), .O(n4406) );
  AOI22S U5595 ( .A1(window_1__4__5_), .A2(n4385), .B1(SRAM_out_buffer[37]), 
        .B2(n4416), .O(n4405) );
  AOI22S U5596 ( .A1(SRAM_out_buffer[45]), .A2(n4709), .B1(SRAM_out_buffer[77]), .B2(n4708), .O(n4404) );
  ND2S U5597 ( .I1(SRAM_out_buffer[68]), .I2(n4466), .O(n4409) );
  AOI22S U5598 ( .A1(window_1__4__4_), .A2(n4385), .B1(SRAM_out_buffer[36]), 
        .B2(n4416), .O(n4408) );
  AOI22S U5599 ( .A1(SRAM_out_buffer[44]), .A2(n4709), .B1(SRAM_out_buffer[76]), .B2(n4708), .O(n4407) );
  ND2S U5600 ( .I1(SRAM_out_buffer[67]), .I2(n4466), .O(n4412) );
  AOI22S U5601 ( .A1(window_1__4__3_), .A2(n4385), .B1(SRAM_out_buffer[35]), 
        .B2(n4416), .O(n4411) );
  AOI22S U5602 ( .A1(SRAM_out_buffer[43]), .A2(n4709), .B1(SRAM_out_buffer[75]), .B2(n4708), .O(n4410) );
  ND2S U5603 ( .I1(SRAM_out_buffer[70]), .I2(n4466), .O(n4415) );
  AOI22S U5604 ( .A1(window_1__4__6_), .A2(n4385), .B1(SRAM_out_buffer[38]), 
        .B2(n4416), .O(n4414) );
  AOI22S U5605 ( .A1(SRAM_out_buffer[46]), .A2(n4709), .B1(SRAM_out_buffer[78]), .B2(n4698), .O(n4413) );
  ND2S U5606 ( .I1(SRAM_out_buffer[71]), .I2(n4466), .O(n4419) );
  AOI22S U5607 ( .A1(window_1__4__7_), .A2(n4385), .B1(SRAM_out_buffer[39]), 
        .B2(n4416), .O(n4418) );
  AOI22S U5608 ( .A1(SRAM_out_buffer[47]), .A2(n4709), .B1(SRAM_out_buffer[79]), .B2(n4698), .O(n4417) );
  AOI22S U5609 ( .A1(n4193), .A2(SRAM_64X32_out_decode[5]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[29]), .O(n4421) );
  AOI22S U5610 ( .A1(n3485), .A2(SRAM_192X32_out_decode[5]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[29]), .O(n4420) );
  MOAI1 U5611 ( .A1(n5675), .A2(n4422), .B1(n5675), .B2(n4422), .O(n6047) );
  INV1S U5612 ( .I(n6047), .O(n5950) );
  AOI22S U5613 ( .A1(n5950), .A2(n4749), .B1(SRAM_out_buffer[29]), .B2(n4771), 
        .O(n5917) );
  AOI22S U5614 ( .A1(median_in[5]), .A2(n4981), .B1(median_in[13]), .B2(n6064), 
        .O(n4423) );
  AOI22S U5615 ( .A1(n4743), .A2(SRAM_192X32_out_decode[30]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[30]), .O(n4425) );
  AOI22S U5616 ( .A1(n4193), .A2(SRAM_64X32_out_decode[6]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[6]), .O(n4424) );
  MOAI1S U5617 ( .A1(n4748), .A2(n4426), .B1(n4746), .B2(n4426), .O(n5967) );
  AOI22S U5618 ( .A1(n5967), .A2(n4749), .B1(SRAM_out_buffer[30]), .B2(n4771), 
        .O(n4437) );
  AOI22S U5619 ( .A1(median_in[14]), .A2(n6064), .B1(median_in[6]), .B2(n4981), 
        .O(n4427) );
  AOI22S U5620 ( .A1(n3485), .A2(SRAM_192X32_out_decode[2]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[26]), .O(n4429) );
  AOI22S U5621 ( .A1(n4193), .A2(SRAM_64X32_out_decode[2]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[26]), .O(n4428) );
  ND2S U5622 ( .I1(n4429), .I2(n4428), .O(n4430) );
  MOAI1 U5623 ( .A1(n4748), .A2(n4430), .B1(n4748), .B2(n4430), .O(n5961) );
  AOI22S U5624 ( .A1(n5961), .A2(n4749), .B1(SRAM_out_buffer[26]), .B2(n4771), 
        .O(n4441) );
  AOI22S U5625 ( .A1(median_in[10]), .A2(n6064), .B1(median_in[2]), .B2(n4981), 
        .O(n4431) );
  INV1S U5626 ( .I(n6037), .O(n5886) );
  AOI22S U5627 ( .A1(window_2__3__2_), .A2(n4889), .B1(n5886), .B2(n4749), .O(
        n4436) );
  INV1S U5628 ( .I(SRAM_out_buffer[58]), .O(n4937) );
  AOI22S U5629 ( .A1(median_in[2]), .A2(n6064), .B1(n4776), .B2(
        SRAM_out_buffer[50]), .O(n4433) );
  OA12S U5630 ( .B1(n4688), .B2(n4937), .A1(n4433), .O(n4435) );
  INV1S U5631 ( .I(n4773), .O(n4751) );
  AOI22S U5632 ( .A1(SRAM_out_buffer[18]), .A2(n4771), .B1(n4751), .B2(n5961), 
        .O(n4434) );
  ND2S U5633 ( .I1(median_in[22]), .I2(n6064), .O(n4440) );
  INV1S U5634 ( .I(n4981), .O(n6068) );
  ND2S U5635 ( .I1(median_in[18]), .I2(n6064), .O(n4444) );
  AOI22S U5636 ( .A1(n4743), .A2(SRAM_192X32_out_decode[25]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[25]), .O(n4446) );
  AOI22S U5637 ( .A1(n4193), .A2(SRAM_64X32_out_decode[1]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[1]), .O(n4445) );
  ND2S U5638 ( .I1(n4446), .I2(n4445), .O(n4447) );
  MOAI1 U5639 ( .A1(n5675), .A2(n4447), .B1(n5675), .B2(n4447), .O(n6035) );
  INV1S U5640 ( .I(n4749), .O(n4892) );
  INV1S U5641 ( .I(SRAM_out_buffer[25]), .O(n5888) );
  INV1S U5642 ( .I(n4448), .O(n4893) );
  OAI22S U5643 ( .A1(n6035), .A2(n4892), .B1(n5888), .B2(n4893), .O(n4978) );
  AOI22S U5644 ( .A1(median_in[9]), .A2(n6064), .B1(median_in[1]), .B2(n4981), 
        .O(n4449) );
  AOI22S U5645 ( .A1(n3485), .A2(SRAM_192X32_out_decode[7]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[31]), .O(n4451) );
  AOI22S U5646 ( .A1(n4193), .A2(SRAM_64X32_out_decode[7]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[31]), .O(n4450) );
  MOAI1 U5647 ( .A1(n5675), .A2(n4452), .B1(n5675), .B2(n4452), .O(n6059) );
  INV1S U5648 ( .I(SRAM_out_buffer[31]), .O(n6058) );
  OAI22S U5649 ( .A1(n6059), .A2(n4892), .B1(n6058), .B2(n4893), .O(n6063) );
  AOI22S U5650 ( .A1(median_in[15]), .A2(n6064), .B1(median_in[7]), .B2(n4981), 
        .O(n4453) );
  INV1S U5651 ( .I(n4455), .O(n61300) );
  AOI22S U5652 ( .A1(SRAM_out_buffer[62]), .A2(n4772), .B1(n4751), .B2(n5967), 
        .O(n4462) );
  MOAI1S U5653 ( .A1(n5942), .A2(n6322), .B1(n4767), .B2(SRAM_out_buffer[54]), 
        .O(n4456) );
  OAI22S U5654 ( .A1(n4889), .A2(n4456), .B1(window_2__3__6_), .B2(n4456), .O(
        n4461) );
  AOI22S U5655 ( .A1(n3485), .A2(SRAM_192X32_out_decode[14]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[22]), .O(n4458) );
  AOI22S U5656 ( .A1(n4193), .A2(SRAM_64X32_out_decode[14]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[22]), .O(n4457) );
  MOAI1 U5657 ( .A1(n5675), .A2(n4459), .B1(n5675), .B2(n4459), .O(n6049) );
  INV1S U5658 ( .I(n6049), .O(n5949) );
  AOI22S U5659 ( .A1(SRAM_out_buffer[22]), .A2(n4771), .B1(n5949), .B2(n4749), 
        .O(n4460) );
  AOI22S U5660 ( .A1(n4193), .A2(SRAM_64X32_out_decode[24]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[0]), .O(n4464) );
  AOI22S U5661 ( .A1(n3485), .A2(SRAM_192X32_out_decode[24]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[0]), .O(n4463) );
  INV1S U5662 ( .I(n5861), .O(n5765) );
  AOI22S U5663 ( .A1(SRAM_out_buffer[40]), .A2(n4772), .B1(n5765), .B2(n4749), 
        .O(n4469) );
  AOI22S U5664 ( .A1(window_2__4__0_), .A2(n4385), .B1(n4751), .B2(n5805), .O(
        n4468) );
  AOI22S U5665 ( .A1(SRAM_out_buffer[0]), .A2(n5770), .B1(SRAM_out_buffer[32]), 
        .B2(n4504), .O(n4467) );
  AOI22S U5666 ( .A1(n4743), .A2(SRAM_192X32_out_decode[7]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[7]), .O(n4471) );
  AOI22S U5667 ( .A1(n4193), .A2(SRAM_64X32_out_decode[31]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[31]), .O(n4470) );
  MOAI1S U5668 ( .A1(n4748), .A2(n4472), .B1(n4746), .B2(n4472), .O(n5850) );
  AOI22S U5669 ( .A1(SRAM_out_buffer[47]), .A2(n4772), .B1(n5850), .B2(n4749), 
        .O(n4475) );
  INV1S U5670 ( .I(n5857), .O(n5884) );
  AOI22S U5671 ( .A1(SRAM_out_buffer[7]), .A2(n5770), .B1(n4751), .B2(n5884), 
        .O(n4474) );
  AOI22S U5672 ( .A1(SRAM_out_buffer[39]), .A2(n4504), .B1(window_2__4__7_), 
        .B2(n4385), .O(n4473) );
  AOI22S U5673 ( .A1(SRAM_out_buffer[42]), .A2(n4772), .B1(n5806), .B2(n4749), 
        .O(n4478) );
  INV1S U5674 ( .I(n5866), .O(n5800) );
  AOI22S U5675 ( .A1(window_2__4__2_), .A2(n4385), .B1(n4751), .B2(n5800), .O(
        n4477) );
  AOI22S U5676 ( .A1(SRAM_out_buffer[2]), .A2(n5770), .B1(SRAM_out_buffer[34]), 
        .B2(n4504), .O(n4476) );
  AOI22S U5677 ( .A1(n3485), .A2(SRAM_192X32_out_decode[28]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[4]), .O(n4480) );
  AOI22S U5678 ( .A1(n4193), .A2(SRAM_64X32_out_decode[28]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[4]), .O(n4479) );
  MOAI1S U5679 ( .A1(n4746), .A2(n4481), .B1(n4748), .B2(n4481), .O(n5793) );
  AOI22S U5680 ( .A1(SRAM_out_buffer[44]), .A2(n4772), .B1(n5793), .B2(n4749), 
        .O(n4487) );
  AOI22S U5681 ( .A1(n4743), .A2(SRAM_192X32_out_decode[12]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[12]), .O(n4483) );
  AOI22S U5682 ( .A1(n4193), .A2(SRAM_64X32_out_decode[20]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[20]), .O(n4482) );
  MOAI1 U5683 ( .A1(n5675), .A2(n4484), .B1(n5675), .B2(n4484), .O(n5872) );
  INV1S U5684 ( .I(n5872), .O(n5798) );
  AOI22S U5685 ( .A1(SRAM_out_buffer[4]), .A2(n5770), .B1(n4751), .B2(n5798), 
        .O(n4486) );
  AOI22S U5686 ( .A1(SRAM_out_buffer[36]), .A2(n4504), .B1(window_2__4__4_), 
        .B2(n4385), .O(n4485) );
  AOI22S U5687 ( .A1(SRAM_out_buffer[46]), .A2(n4772), .B1(n5813), .B2(n4749), 
        .O(n4490) );
  INV1S U5688 ( .I(n5878), .O(n5772) );
  AOI22S U5689 ( .A1(SRAM_out_buffer[6]), .A2(n5770), .B1(n4751), .B2(n5772), 
        .O(n4489) );
  AOI22S U5690 ( .A1(SRAM_out_buffer[38]), .A2(n4504), .B1(window_2__4__6_), 
        .B2(n4385), .O(n4488) );
  INV1S U5691 ( .I(n5869), .O(n5797) );
  AOI22S U5692 ( .A1(SRAM_out_buffer[43]), .A2(n4772), .B1(n4751), .B2(n5797), 
        .O(n4493) );
  AOI22S U5693 ( .A1(SRAM_out_buffer[3]), .A2(n5770), .B1(n5799), .B2(n4749), 
        .O(n4492) );
  AOI22S U5694 ( .A1(SRAM_out_buffer[35]), .A2(n4504), .B1(window_2__4__3_), 
        .B2(n4385), .O(n4491) );
  AOI22S U5695 ( .A1(SRAM_out_buffer[45]), .A2(n4772), .B1(n5791), .B2(n4749), 
        .O(n4496) );
  INV1S U5696 ( .I(n5875), .O(n5792) );
  AOI22S U5697 ( .A1(window_2__4__5_), .A2(n4385), .B1(n4751), .B2(n5792), .O(
        n4495) );
  AOI22S U5698 ( .A1(SRAM_out_buffer[5]), .A2(n5770), .B1(SRAM_out_buffer[37]), 
        .B2(n4504), .O(n4494) );
  AOI22S U5699 ( .A1(SRAM_out_buffer[56]), .A2(n4772), .B1(n4751), .B2(n5964), 
        .O(n4503) );
  INV1S U5700 ( .I(median_in[0]), .O(n5262) );
  MOAI1S U5701 ( .A1(n5942), .A2(n5262), .B1(n4767), .B2(SRAM_out_buffer[48]), 
        .O(n4497) );
  OAI22S U5702 ( .A1(n4889), .A2(n4497), .B1(window_2__3__0_), .B2(n4497), .O(
        n4502) );
  AOI22S U5703 ( .A1(n4193), .A2(SRAM_64X32_out_decode[8]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[16]), .O(n4499) );
  AOI22S U5704 ( .A1(n3485), .A2(SRAM_192X32_out_decode[8]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[16]), .O(n4498) );
  ND2S U5705 ( .I1(n4499), .I2(n4498), .O(n4500) );
  MOAI1 U5706 ( .A1(n5675), .A2(n4500), .B1(n5675), .B2(n4500), .O(n6031) );
  INV1S U5707 ( .I(n6031), .O(n5885) );
  AOI22S U5708 ( .A1(SRAM_out_buffer[16]), .A2(n4771), .B1(n5885), .B2(n4749), 
        .O(n4501) );
  INV1S U5709 ( .I(n5864), .O(n5807) );
  AOI22S U5710 ( .A1(SRAM_out_buffer[41]), .A2(n4772), .B1(n5807), .B2(n4749), 
        .O(n4507) );
  AOI22S U5711 ( .A1(window_2__4__1_), .A2(n4385), .B1(n4751), .B2(n5804), .O(
        n4506) );
  AOI22S U5712 ( .A1(SRAM_out_buffer[1]), .A2(n5770), .B1(SRAM_out_buffer[33]), 
        .B2(n4504), .O(n4505) );
  INV1S U5713 ( .I(n4857), .O(n4508) );
  AOI22S U5714 ( .A1(n4509), .A2(n5767), .B1(n4508), .B2(n3517), .O(n4511) );
  ND2 U5715 ( .I1(n4511), .I2(n4510), .O(n5771) );
  NR2 U5716 ( .I1(n4623), .I2(n4929), .O(n4971) );
  NR2 U5717 ( .I1(n4971), .I2(n4648), .O(n5769) );
  AOI22S U5718 ( .A1(SRAM_out_buffer[88]), .A2(n5771), .B1(SRAM_out_buffer[80]), .B2(n4935), .O(n4515) );
  ND2S U5719 ( .I1(median_in[48]), .I2(n6064), .O(n4513) );
  AOI22S U5720 ( .A1(SRAM_out_buffer[90]), .A2(n5771), .B1(SRAM_out_buffer[82]), .B2(n4935), .O(n4518) );
  ND2S U5721 ( .I1(median_in[50]), .I2(n6064), .O(n4516) );
  AOI22S U5722 ( .A1(n4193), .A2(SRAM_64X32_out_decode[9]), .B1(
        SRAM_192X32_out_decode[17]), .B2(n4743), .O(n4520) );
  AOI22S U5723 ( .A1(SRAM_64X32_out_decode[17]), .A2(n4742), .B1(n3485), .B2(
        SRAM_192X32_out_decode[9]), .O(n4519) );
  ND2S U5724 ( .I1(n4520), .I2(n4519), .O(n4521) );
  MOAI1 U5725 ( .A1(n5675), .A2(n4521), .B1(n5675), .B2(n4521), .O(n6034) );
  MOAI1S U5726 ( .A1(n6034), .A2(n4892), .B1(SRAM_out_buffer[17]), .B2(n4771), 
        .O(n4523) );
  INV1S U5727 ( .I(SRAM_out_buffer[57]), .O(n5889) );
  OAI22S U5728 ( .A1(n6035), .A2(n4773), .B1(n5889), .B2(n4688), .O(n4522) );
  NR2 U5729 ( .I1(n4523), .I2(n4522), .O(n4526) );
  AOI22S U5730 ( .A1(median_in[1]), .A2(n6064), .B1(n4776), .B2(
        SRAM_out_buffer[49]), .O(n4525) );
  NR2 U5731 ( .I1(n5695), .I2(n4547), .O(n4611) );
  ND2P U5732 ( .I1(n3537), .I2(n4611), .O(n4627) );
  NR2 U5733 ( .I1(n3486), .I2(n4627), .O(n4625) );
  INV1S U5734 ( .I(n4527), .O(n4528) );
  INV1S U5735 ( .I(n4529), .O(n4530) );
  NR2 U5736 ( .I1(n4531), .I2(n4547), .O(n4566) );
  AOI22S U5737 ( .A1(n4566), .A2(n6016), .B1(n4620), .B2(n4532), .O(n4533) );
  OAI12HS U5738 ( .B1(n4602), .B2(n4943), .A1(n4533), .O(n4583) );
  INV1S U5739 ( .I(n4583), .O(n4538) );
  AOI22S U5740 ( .A1(n5985), .A2(n4566), .B1(n4620), .B2(n4550), .O(n4575) );
  INV1S U5741 ( .I(n4620), .O(n4617) );
  NR2 U5742 ( .I1(n4535), .I2(n4617), .O(n4536) );
  NR2 U5743 ( .I1(n4587), .I2(n4536), .O(n4537) );
  NR2 U5744 ( .I1(n4540), .I2(n4562), .O(n4580) );
  ND3S U5745 ( .I1(n4542), .I2(n5766), .I3(n4541), .O(n4574) );
  ND3P U5746 ( .I1(n4543), .I2(n4552), .I3(n4574), .O(n5122) );
  XOR2HS U5747 ( .I1(n4544), .I2(n5122), .O(n4737) );
  NR2 U5748 ( .I1(n4548), .I2(n4547), .O(n4565) );
  AOI22S U5749 ( .A1(n5985), .A2(n4565), .B1(n4620), .B2(n4549), .O(n4551) );
  ND2S U5750 ( .I1(n4625), .I2(n4550), .O(n4594) );
  AN4B1S U5751 ( .I1(n4552), .I2(n4551), .I3(n4594), .B1(n4587), .O(n4576) );
  NR2 U5752 ( .I1(n4553), .I2(n4627), .O(n4612) );
  ND2S U5753 ( .I1(n4612), .I2(n4554), .O(n4559) );
  AOI22S U5754 ( .A1(n6016), .A2(n4565), .B1(n4625), .B2(n4555), .O(n4558) );
  ND2S U5755 ( .I1(n4620), .I2(n4556), .O(n4557) );
  ND3S U5756 ( .I1(n4559), .I2(n4558), .I3(n4557), .O(n4586) );
  NR2 U5757 ( .I1(n4580), .I2(n4586), .O(n4560) );
  ND2S U5758 ( .I1(n4576), .I2(n4560), .O(n4561) );
  XOR2HS U5759 ( .I1(n4561), .I2(n5122), .O(n5108) );
  ND2S U5760 ( .I1(n5766), .I2(n4564), .O(n4567) );
  MOAI1S U5761 ( .A1(n4627), .A2(n4567), .B1(n4630), .B2(n5743), .O(n4568) );
  AOI12HS U5762 ( .B1(n4625), .B2(n4569), .A1(n4568), .O(n4572) );
  ND2S U5763 ( .I1(n4612), .I2(n4570), .O(n4571) );
  ND3S U5764 ( .I1(n4573), .I2(n4572), .I3(n4571), .O(n4579) );
  INV1S U5765 ( .I(n4574), .O(n4592) );
  AN3B2S U5766 ( .I1(n4575), .B1(n4579), .B2(n4592), .O(n4577) );
  ND2S U5767 ( .I1(n4577), .I2(n4576), .O(n4578) );
  XOR2HS U5768 ( .I1(n4578), .I2(n5122), .O(n5121) );
  NR2 U5769 ( .I1(n4580), .I2(n4579), .O(n4590) );
  NR2 U5770 ( .I1(n4584), .I2(n4583), .O(n4589) );
  NR2 U5771 ( .I1(n4585), .I2(n4617), .O(n4735) );
  NR3 U5772 ( .I1(n4587), .I2(n4735), .I3(n4586), .O(n4588) );
  NR2 U5773 ( .I1(n4592), .I2(n4591), .O(n4595) );
  OAI112HS U5774 ( .C1(n4599), .C2(n4627), .A1(n4598), .B1(n4597), .O(n4600)
         );
  NR2 U5775 ( .I1(n4601), .I2(n4600), .O(n5126) );
  INV1S U5776 ( .I(n4602), .O(n4603) );
  OAI12HS U5777 ( .B1(n4605), .B2(n4604), .A1(n4603), .O(n4616) );
  OA13S U5778 ( .B1(n4618), .B2(n4617), .B3(n4606), .A1(n4616), .O(n4607) );
  MOAI1S U5779 ( .A1(n4608), .A2(n4607), .B1(n6015), .B2(n4630), .O(n4609) );
  AOI13HS U5780 ( .B1(n5918), .B2(n4611), .B3(n4610), .A1(n4609), .O(n4615) );
  OAI112HS U5781 ( .C1(n6245), .C2(n4613), .A1(n4612), .B1(n5727), .O(n4614)
         );
  AOI22S U5782 ( .A1(n5126), .A2(SRAM_64X32_addr[2]), .B1(n5124), .B2(N1045), 
        .O(n4635) );
  MOAI1S U5783 ( .A1(n4622), .A2(n4621), .B1(n4620), .B2(n4619), .O(n4629) );
  INV1S U5784 ( .I(n5721), .O(n4626) );
  INV1S U5785 ( .I(n4623), .O(n4624) );
  MOAI1S U5786 ( .A1(n4627), .A2(n4626), .B1(n4625), .B2(n4624), .O(n4628) );
  NR2 U5787 ( .I1(n4629), .I2(n4628), .O(n4633) );
  AOI22S U5788 ( .A1(n3485), .A2(SRAM_192X32_out_decode[11]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[19]), .O(n4638) );
  AOI22S U5789 ( .A1(n4193), .A2(SRAM_64X32_out_decode[11]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[19]), .O(n4637) );
  MOAI1 U5790 ( .A1(n5675), .A2(n4639), .B1(n5675), .B2(n4639), .O(n6040) );
  INV1S U5791 ( .I(n6040), .O(n5887) );
  AOI22S U5792 ( .A1(window_2__3__3_), .A2(n4889), .B1(n5887), .B2(n4749), .O(
        n4646) );
  INV1S U5793 ( .I(SRAM_out_buffer[59]), .O(n5898) );
  MOAI1S U5794 ( .A1(n5898), .A2(n4688), .B1(n6064), .B2(median_in[3]), .O(
        n4640) );
  OAI22S U5795 ( .A1(n4776), .A2(n4640), .B1(SRAM_out_buffer[51]), .B2(n4640), 
        .O(n4645) );
  AOI22S U5796 ( .A1(n4193), .A2(SRAM_64X32_out_decode[3]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[27]), .O(n4642) );
  AOI22S U5797 ( .A1(n3485), .A2(SRAM_192X32_out_decode[3]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[27]), .O(n4641) );
  ND2S U5798 ( .I1(n4642), .I2(n4641), .O(n4643) );
  MOAI1S U5799 ( .A1(n4748), .A2(n4643), .B1(n4748), .B2(n4643), .O(n5956) );
  AOI22S U5800 ( .A1(SRAM_out_buffer[19]), .A2(n4771), .B1(n4751), .B2(n5956), 
        .O(n4644) );
  AOI22S U5801 ( .A1(median_in[27]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[83]), .O(n4651) );
  AOI22S U5802 ( .A1(n4709), .A2(SRAM_out_buffer[59]), .B1(SRAM_out_buffer[91]), .B2(n4708), .O(n4650) );
  NR2 U5803 ( .I1(n4771), .I2(n4648), .O(n4938) );
  AOI22S U5804 ( .A1(window_1__3__3_), .A2(n4889), .B1(SRAM_out_buffer[51]), 
        .B2(n4914), .O(n4649) );
  AOI22S U5805 ( .A1(median_in[28]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[84]), .O(n4654) );
  AOI22S U5806 ( .A1(n4709), .A2(SRAM_out_buffer[60]), .B1(SRAM_out_buffer[92]), .B2(n4708), .O(n4653) );
  AOI22S U5807 ( .A1(window_1__3__4_), .A2(n4889), .B1(SRAM_out_buffer[52]), 
        .B2(n4914), .O(n4652) );
  AOI22S U5808 ( .A1(median_in[30]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[86]), .O(n4657) );
  AOI22S U5809 ( .A1(n4709), .A2(SRAM_out_buffer[62]), .B1(SRAM_out_buffer[94]), .B2(n4708), .O(n4656) );
  AOI22S U5810 ( .A1(window_1__3__6_), .A2(n4889), .B1(SRAM_out_buffer[54]), 
        .B2(n4914), .O(n4655) );
  AOI22S U5811 ( .A1(median_in[31]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[87]), .O(n4660) );
  AOI22S U5812 ( .A1(n4709), .A2(SRAM_out_buffer[63]), .B1(SRAM_out_buffer[95]), .B2(n4708), .O(n4659) );
  AOI22S U5813 ( .A1(window_1__3__7_), .A2(n4889), .B1(SRAM_out_buffer[55]), 
        .B2(n4914), .O(n4658) );
  AOI22S U5814 ( .A1(SRAM_out_buffer[79]), .A2(n5935), .B1(window_1__3__7_), 
        .B2(n6064), .O(n4663) );
  AOI22S U5815 ( .A1(SRAM_out_buffer[55]), .A2(n4709), .B1(SRAM_out_buffer[87]), .B2(n4708), .O(n4662) );
  AOI22S U5816 ( .A1(window_1__4__7_), .A2(n4889), .B1(SRAM_out_buffer[47]), 
        .B2(n4914), .O(n4661) );
  AOI22S U5817 ( .A1(SRAM_out_buffer[75]), .A2(n5935), .B1(window_1__3__3_), 
        .B2(n6064), .O(n4666) );
  AOI22S U5818 ( .A1(SRAM_out_buffer[51]), .A2(n4709), .B1(SRAM_out_buffer[83]), .B2(n4698), .O(n4665) );
  AOI22S U5819 ( .A1(window_1__4__3_), .A2(n4889), .B1(SRAM_out_buffer[43]), 
        .B2(n4914), .O(n4664) );
  AOI22S U5820 ( .A1(SRAM_out_buffer[73]), .A2(n5935), .B1(window_1__3__1_), 
        .B2(n6064), .O(n4669) );
  AOI22S U5821 ( .A1(SRAM_out_buffer[49]), .A2(n4709), .B1(SRAM_out_buffer[81]), .B2(n4708), .O(n4668) );
  AOI22S U5822 ( .A1(window_1__4__1_), .A2(n4889), .B1(SRAM_out_buffer[41]), 
        .B2(n4914), .O(n4667) );
  AOI22S U5823 ( .A1(SRAM_out_buffer[76]), .A2(n5935), .B1(window_1__3__4_), 
        .B2(n6064), .O(n4672) );
  AOI22S U5824 ( .A1(SRAM_out_buffer[52]), .A2(n4709), .B1(SRAM_out_buffer[84]), .B2(n4698), .O(n4671) );
  AOI22S U5825 ( .A1(window_1__4__4_), .A2(n4889), .B1(SRAM_out_buffer[44]), 
        .B2(n4914), .O(n4670) );
  AOI22S U5826 ( .A1(SRAM_out_buffer[77]), .A2(n5935), .B1(window_1__3__5_), 
        .B2(n6064), .O(n4675) );
  AOI22S U5827 ( .A1(SRAM_out_buffer[53]), .A2(n4709), .B1(SRAM_out_buffer[85]), .B2(n4708), .O(n4674) );
  AOI22S U5828 ( .A1(window_1__4__5_), .A2(n4889), .B1(SRAM_out_buffer[45]), 
        .B2(n4914), .O(n4673) );
  AOI22S U5829 ( .A1(SRAM_out_buffer[74]), .A2(n5935), .B1(window_1__3__2_), 
        .B2(n6064), .O(n4678) );
  AOI22S U5830 ( .A1(SRAM_out_buffer[50]), .A2(n4709), .B1(SRAM_out_buffer[82]), .B2(n4698), .O(n4677) );
  AOI22S U5831 ( .A1(window_1__4__2_), .A2(n4889), .B1(SRAM_out_buffer[42]), 
        .B2(n4914), .O(n4676) );
  AOI22S U5832 ( .A1(SRAM_out_buffer[78]), .A2(n5935), .B1(window_1__3__6_), 
        .B2(n6064), .O(n4681) );
  AOI22S U5833 ( .A1(SRAM_out_buffer[54]), .A2(n4709), .B1(SRAM_out_buffer[86]), .B2(n4708), .O(n4680) );
  AOI22S U5834 ( .A1(window_1__4__6_), .A2(n4889), .B1(SRAM_out_buffer[46]), 
        .B2(n4914), .O(n4679) );
  MOAI1S U5835 ( .A1(n6059), .A2(n4773), .B1(SRAM_out_buffer[23]), .B2(n4771), 
        .O(n4683) );
  NR2 U5836 ( .I1(n5942), .I2(n5276), .O(n4682) );
  NR2 U5837 ( .I1(n4683), .I2(n4682), .O(n4686) );
  AOI22S U5838 ( .A1(SRAM_out_buffer[63]), .A2(n4772), .B1(n5969), .B2(n4749), 
        .O(n4685) );
  AOI22S U5839 ( .A1(n4776), .A2(SRAM_out_buffer[55]), .B1(n4889), .B2(
        window_2__3__7_), .O(n4684) );
  AOI22S U5840 ( .A1(window_2__3__4_), .A2(n4889), .B1(n4751), .B2(n5955), .O(
        n4694) );
  INV1S U5841 ( .I(SRAM_out_buffer[60]), .O(n4861) );
  AOI22S U5842 ( .A1(median_in[4]), .A2(n6064), .B1(n4776), .B2(
        SRAM_out_buffer[52]), .O(n4687) );
  OA12S U5843 ( .B1(n4688), .B2(n4861), .A1(n4687), .O(n4693) );
  AOI22S U5844 ( .A1(n3485), .A2(SRAM_192X32_out_decode[12]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[20]), .O(n4690) );
  AOI22S U5845 ( .A1(n4193), .A2(SRAM_64X32_out_decode[12]), .B1(n4743), .B2(
        SRAM_192X32_out_decode[20]), .O(n4689) );
  MOAI1S U5846 ( .A1(n4746), .A2(n4691), .B1(n4746), .B2(n4691), .O(n5951) );
  AOI22S U5847 ( .A1(SRAM_out_buffer[20]), .A2(n4771), .B1(n5951), .B2(n4749), 
        .O(n4692) );
  AOI22S U5848 ( .A1(window_1__3__2_), .A2(n4889), .B1(SRAM_out_buffer[50]), 
        .B2(n4914), .O(n4697) );
  AOI22S U5849 ( .A1(n4709), .A2(SRAM_out_buffer[58]), .B1(SRAM_out_buffer[90]), .B2(n4708), .O(n4696) );
  AOI22S U5850 ( .A1(n6064), .A2(median_in[26]), .B1(n5935), .B2(
        SRAM_out_buffer[82]), .O(n4695) );
  AOI22S U5851 ( .A1(window_1__3__1_), .A2(n4889), .B1(SRAM_out_buffer[49]), 
        .B2(n4914), .O(n4701) );
  AOI22S U5852 ( .A1(n4709), .A2(SRAM_out_buffer[57]), .B1(SRAM_out_buffer[89]), .B2(n4698), .O(n4700) );
  AOI22S U5853 ( .A1(median_in[25]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[81]), .O(n4699) );
  AOI22S U5854 ( .A1(window_1__3__0_), .A2(n4889), .B1(SRAM_out_buffer[48]), 
        .B2(n4914), .O(n4704) );
  AOI22S U5855 ( .A1(SRAM_out_buffer[88]), .A2(n4708), .B1(SRAM_out_buffer[56]), .B2(n4709), .O(n4703) );
  AOI22S U5856 ( .A1(median_in[24]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[80]), .O(n4702) );
  AOI22S U5857 ( .A1(SRAM_out_buffer[72]), .A2(n5935), .B1(window_1__3__0_), 
        .B2(n6064), .O(n4707) );
  AOI22S U5858 ( .A1(n4709), .A2(SRAM_out_buffer[48]), .B1(SRAM_out_buffer[80]), .B2(n4708), .O(n4706) );
  AOI22S U5859 ( .A1(window_1__4__0_), .A2(n4889), .B1(SRAM_out_buffer[40]), 
        .B2(n4914), .O(n4705) );
  AOI22S U5860 ( .A1(median_in[29]), .A2(n6064), .B1(n5935), .B2(
        SRAM_out_buffer[85]), .O(n4712) );
  AOI22S U5861 ( .A1(n4709), .A2(SRAM_out_buffer[61]), .B1(SRAM_out_buffer[93]), .B2(n4708), .O(n4711) );
  AOI22S U5862 ( .A1(window_1__3__5_), .A2(n4889), .B1(SRAM_out_buffer[53]), 
        .B2(n4914), .O(n4710) );
  HA1 U5863 ( .A(conv_temp[17]), .B(n4713), .C(n4780), .S(n4714) );
  INV1S U5864 ( .I(n4714), .O(n61290) );
  MOAI1S U5865 ( .A1(n6031), .A2(n4773), .B1(SRAM_out_buffer[8]), .B2(n4771), 
        .O(n4716) );
  MOAI1S U5866 ( .A1(n5860), .A2(n4892), .B1(window_2__4__0_), .B2(n4889), .O(
        n4715) );
  NR2 U5867 ( .I1(n4716), .I2(n4715), .O(n4719) );
  AOI22S U5868 ( .A1(SRAM_out_buffer[40]), .A2(n4776), .B1(window_2__3__0_), 
        .B2(n6064), .O(n4718) );
  MOAI1S U5869 ( .A1(n6037), .A2(n4773), .B1(SRAM_out_buffer[10]), .B2(n4771), 
        .O(n4721) );
  MOAI1S U5870 ( .A1(n5866), .A2(n4892), .B1(window_2__4__2_), .B2(n4889), .O(
        n4720) );
  NR2 U5871 ( .I1(n4721), .I2(n4720), .O(n4724) );
  AOI22S U5872 ( .A1(SRAM_out_buffer[50]), .A2(n4772), .B1(window_2__3__2_), 
        .B2(n6064), .O(n4723) );
  MOAI1S U5873 ( .A1(n6049), .A2(n4773), .B1(SRAM_out_buffer[14]), .B2(n4771), 
        .O(n4726) );
  MOAI1S U5874 ( .A1(n5878), .A2(n4892), .B1(window_2__4__6_), .B2(n4889), .O(
        n4725) );
  NR2 U5875 ( .I1(n4726), .I2(n4725), .O(n4729) );
  AOI22S U5876 ( .A1(n4776), .A2(SRAM_out_buffer[46]), .B1(SRAM_out_buffer[54]), .B2(n4772), .O(n4728) );
  ND2S U5877 ( .I1(window_2__3__6_), .I2(n6064), .O(n4727) );
  MOAI1S U5878 ( .A1(n5857), .A2(n4892), .B1(SRAM_out_buffer[15]), .B2(n4771), 
        .O(n4731) );
  MOAI1S U5879 ( .A1(n6029), .A2(n4773), .B1(window_2__4__7_), .B2(n4889), .O(
        n4730) );
  NR2 U5880 ( .I1(n4731), .I2(n4730), .O(n4734) );
  AOI22S U5881 ( .A1(SRAM_out_buffer[47]), .A2(n4776), .B1(window_2__3__7_), 
        .B2(n6064), .O(n4733) );
  XOR2HS U5882 ( .I1(n4735), .I2(n5122), .O(n4923) );
  FA1 U5883 ( .A(N1045), .B(n4737), .CI(n4736), .CO(n4922), .S(n4596) );
  AOI22S U5884 ( .A1(n5126), .A2(SRAM_64X32_addr[3]), .B1(n5124), .B2(N1046), 
        .O(n4740) );
  AOI22S U5885 ( .A1(n4193), .A2(SRAM_64X32_out_decode[13]), .B1(n3485), .B2(
        SRAM_192X32_out_decode[13]), .O(n4745) );
  AOI22S U5886 ( .A1(n4743), .A2(SRAM_192X32_out_decode[21]), .B1(n4742), .B2(
        SRAM_64X32_out_decode[21]), .O(n4744) );
  MOAI1S U5887 ( .A1(n4748), .A2(n4747), .B1(n4746), .B2(n4747), .O(n5948) );
  AOI22S U5888 ( .A1(SRAM_out_buffer[61]), .A2(n4772), .B1(n5948), .B2(n4749), 
        .O(n4754) );
  INV1S U5889 ( .I(median_in[5]), .O(n5269) );
  AOI22S U5890 ( .A1(n4767), .A2(SRAM_out_buffer[53]), .B1(n4889), .B2(
        window_2__3__5_), .O(n4750) );
  AOI22S U5891 ( .A1(SRAM_out_buffer[21]), .A2(n4771), .B1(n4751), .B2(n5950), 
        .O(n4752) );
  MOAI1S U5892 ( .A1(n6034), .A2(n4773), .B1(SRAM_out_buffer[9]), .B2(n4771), 
        .O(n4756) );
  MOAI1S U5893 ( .A1(n5863), .A2(n4892), .B1(SRAM_out_buffer[49]), .B2(n4772), 
        .O(n4755) );
  NR2 U5894 ( .I1(n4756), .I2(n4755), .O(n4759) );
  AOI22S U5895 ( .A1(window_2__4__1_), .A2(n4889), .B1(window_2__3__1_), .B2(
        n6064), .O(n4758) );
  ND2S U5896 ( .I1(n4767), .I2(SRAM_out_buffer[41]), .O(n4757) );
  INV1S U5897 ( .I(n5948), .O(n6046) );
  MOAI1S U5898 ( .A1(n6046), .A2(n4773), .B1(SRAM_out_buffer[13]), .B2(n4771), 
        .O(n4761) );
  MOAI1S U5899 ( .A1(n5875), .A2(n4892), .B1(SRAM_out_buffer[53]), .B2(n4772), 
        .O(n4760) );
  NR2 U5900 ( .I1(n4761), .I2(n4760), .O(n4764) );
  AOI22S U5901 ( .A1(n4776), .A2(SRAM_out_buffer[45]), .B1(n4889), .B2(
        window_2__4__5_), .O(n4763) );
  ND2S U5902 ( .I1(window_2__3__5_), .I2(n6064), .O(n4762) );
  INV1S U5903 ( .I(n5951), .O(n6043) );
  MOAI1S U5904 ( .A1(n6043), .A2(n4773), .B1(SRAM_out_buffer[12]), .B2(n4771), 
        .O(n4766) );
  MOAI1S U5905 ( .A1(n5872), .A2(n4892), .B1(SRAM_out_buffer[52]), .B2(n4772), 
        .O(n4765) );
  NR2 U5906 ( .I1(n4766), .I2(n4765), .O(n4770) );
  AOI22S U5907 ( .A1(window_2__4__4_), .A2(n4889), .B1(window_2__3__4_), .B2(
        n6064), .O(n4769) );
  ND2S U5908 ( .I1(n4767), .I2(SRAM_out_buffer[44]), .O(n4768) );
  MOAI1S U5909 ( .A1(n5869), .A2(n4892), .B1(SRAM_out_buffer[11]), .B2(n4771), 
        .O(n4775) );
  MOAI1S U5910 ( .A1(n6040), .A2(n4773), .B1(SRAM_out_buffer[51]), .B2(n4772), 
        .O(n4774) );
  NR2 U5911 ( .I1(n4775), .I2(n4774), .O(n4779) );
  AOI22S U5912 ( .A1(SRAM_out_buffer[43]), .A2(n4776), .B1(window_2__3__3_), 
        .B2(n6064), .O(n4778) );
  HA1P U5913 ( .A(conv_temp[18]), .B(n4780), .C(n3888), .S(n4781) );
  ND2S U5914 ( .I1(start_write_flag), .I2(n5095), .O(n4783) );
  ND2S U5915 ( .I1(SRAM_192_32_in_count[0]), .I2(SRAM_192_32_in_count[1]), .O(
        n5648) );
  ND2S U5916 ( .I1(n4783), .I2(n5648), .O(n3268) );
  ND2S U5917 ( .I1(n4784), .I2(n5940), .O(find_median_inst_max1[7]) );
  ND2S U5918 ( .I1(n4785), .I2(n5276), .O(find_median_inst_max3[7]) );
  AOI22S U5919 ( .A1(n4854), .A2(gray_avg_reg[5]), .B1(n4799), .B2(
        gray_max_temp[5]), .O(n4790) );
  AOI22S U5920 ( .A1(gray_wgt_reg[5]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[29]), .B2(n4849), .O(n4789) );
  ND2S U5921 ( .I1(n4790), .I2(n4789), .O(n3238) );
  AOI22S U5922 ( .A1(n4854), .A2(gray_avg_reg[4]), .B1(n4799), .B2(
        gray_max_temp[4]), .O(n4792) );
  AOI22S U5923 ( .A1(gray_wgt_reg[4]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[28]), .B2(n4849), .O(n4791) );
  ND2S U5924 ( .I1(n4792), .I2(n4791), .O(n3239) );
  AOI22S U5925 ( .A1(n4854), .A2(gray_avg_reg[6]), .B1(n4799), .B2(
        gray_max_temp[6]), .O(n4794) );
  AOI22S U5926 ( .A1(gray_wgt_reg[6]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[30]), .B2(n4849), .O(n4793) );
  ND2S U5927 ( .I1(n4794), .I2(n4793), .O(n3237) );
  AOI22S U5928 ( .A1(gray_wgt_reg[1]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[25]), .B2(n4849), .O(n4796) );
  AOI22S U5929 ( .A1(n4854), .A2(gray_avg_reg[1]), .B1(n4799), .B2(
        gray_max_temp[1]), .O(n4795) );
  ND2S U5930 ( .I1(n4796), .I2(n4795), .O(n3242) );
  AOI22S U5931 ( .A1(gray_max_temp[29]), .A2(n4799), .B1(gray_avg_reg[29]), 
        .B2(n4854), .O(n4798) );
  AOI22S U5932 ( .A1(gray_wgt_reg[29]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[5]), .B2(n4849), .O(n4797) );
  ND2S U5933 ( .I1(n4798), .I2(n4797), .O(n3262) );
  AOI22S U5934 ( .A1(gray_avg_reg[15]), .A2(n4854), .B1(
        SRAM_192X32_data_in_reg[23]), .B2(n4849), .O(n4801) );
  AOI22S U5935 ( .A1(n4836), .A2(gray_wgt_reg[15]), .B1(n4799), .B2(
        gray_max_temp[15]), .O(n4800) );
  ND2S U5936 ( .I1(n4801), .I2(n4800), .O(n3244) );
  AOI22S U5937 ( .A1(gray_max_temp[31]), .A2(n4799), .B1(
        SRAM_192X32_data_in_reg[7]), .B2(n4849), .O(n4803) );
  AOI22S U5938 ( .A1(n4836), .A2(gray_wgt_reg[31]), .B1(n4854), .B2(
        gray_avg_reg[31]), .O(n4802) );
  ND2S U5939 ( .I1(n4803), .I2(n4802), .O(n3260) );
  AOI22S U5940 ( .A1(n4799), .A2(gray_max_temp[24]), .B1(
        SRAM_192X32_data_in_reg[0]), .B2(n4849), .O(n4805) );
  AOI22S U5941 ( .A1(gray_avg_reg[24]), .A2(n4854), .B1(gray_wgt_reg[24]), 
        .B2(n4836), .O(n4804) );
  ND2S U5942 ( .I1(n4805), .I2(n4804), .O(n3267) );
  AOI22S U5943 ( .A1(n4854), .A2(gray_avg_reg[30]), .B1(
        SRAM_192X32_data_in_reg[6]), .B2(n4849), .O(n4807) );
  AOI22S U5944 ( .A1(gray_max_temp[30]), .A2(n4799), .B1(n4836), .B2(
        gray_wgt_reg[30]), .O(n4806) );
  ND2S U5945 ( .I1(n4807), .I2(n4806), .O(n3261) );
  AOI22S U5946 ( .A1(gray_wgt_reg[27]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[3]), .B2(n4849), .O(n4809) );
  AOI22S U5947 ( .A1(gray_avg_reg[27]), .A2(n4854), .B1(gray_max_temp[27]), 
        .B2(n4799), .O(n4808) );
  ND2S U5948 ( .I1(n4809), .I2(n4808), .O(n3264) );
  AOI22S U5949 ( .A1(gray_wgt_reg[28]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[4]), .B2(n4849), .O(n4811) );
  AOI22S U5950 ( .A1(gray_avg_reg[28]), .A2(n4854), .B1(gray_max_temp[28]), 
        .B2(n4799), .O(n4810) );
  ND2S U5951 ( .I1(n4811), .I2(n4810), .O(n3263) );
  AOI22S U5952 ( .A1(n4836), .A2(gray_wgt_reg[14]), .B1(n4799), .B2(
        gray_max_temp[14]), .O(n4813) );
  AOI22S U5953 ( .A1(gray_avg_reg[14]), .A2(n4854), .B1(
        SRAM_192X32_data_in_reg[22]), .B2(n4849), .O(n4812) );
  ND2S U5954 ( .I1(n4813), .I2(n4812), .O(n3245) );
  AOI22S U5955 ( .A1(gray_avg_reg[25]), .A2(n4854), .B1(n4836), .B2(
        gray_wgt_reg[25]), .O(n4815) );
  AOI22S U5956 ( .A1(n4799), .A2(gray_max_temp[25]), .B1(
        SRAM_192X32_data_in_reg[1]), .B2(n4849), .O(n4814) );
  ND2S U5957 ( .I1(n4815), .I2(n4814), .O(n3266) );
  AOI22S U5958 ( .A1(gray_wgt_reg[17]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[9]), .B2(n4849), .O(n4817) );
  AOI22S U5959 ( .A1(n4854), .A2(gray_avg_reg[17]), .B1(n4799), .B2(
        gray_max_temp[17]), .O(n4816) );
  ND2S U5960 ( .I1(n4817), .I2(n4816), .O(n3258) );
  AOI22S U5961 ( .A1(gray_wgt_reg[22]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[14]), .B2(n4849), .O(n4819) );
  AOI22S U5962 ( .A1(n4854), .A2(gray_avg_reg[22]), .B1(n4799), .B2(
        gray_max_temp[22]), .O(n4818) );
  ND2S U5963 ( .I1(n4819), .I2(n4818), .O(n3253) );
  AOI22S U5964 ( .A1(gray_wgt_reg[19]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[11]), .B2(n4849), .O(n4821) );
  AOI22S U5965 ( .A1(n4854), .A2(gray_avg_reg[19]), .B1(n4799), .B2(
        gray_max_temp[19]), .O(n4820) );
  ND2S U5966 ( .I1(n4821), .I2(n4820), .O(n3256) );
  AOI22S U5967 ( .A1(gray_avg_reg[26]), .A2(n4854), .B1(gray_max_temp[26]), 
        .B2(n4799), .O(n4823) );
  AOI22S U5968 ( .A1(gray_wgt_reg[26]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[2]), .B2(n4849), .O(n4822) );
  ND2S U5969 ( .I1(n4823), .I2(n4822), .O(n3265) );
  AOI22S U5970 ( .A1(n4854), .A2(gray_avg_reg[9]), .B1(n4799), .B2(
        gray_max_temp[9]), .O(n4825) );
  AOI22S U5971 ( .A1(gray_wgt_reg[9]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[17]), .B2(n4849), .O(n4824) );
  ND2S U5972 ( .I1(n4825), .I2(n4824), .O(n3250) );
  AOI22S U5973 ( .A1(n4836), .A2(gray_wgt_reg[13]), .B1(n4799), .B2(
        gray_max_temp[13]), .O(n4827) );
  AOI22S U5974 ( .A1(gray_avg_reg[13]), .A2(n4854), .B1(
        SRAM_192X32_data_in_reg[21]), .B2(n4849), .O(n4826) );
  ND2S U5975 ( .I1(n4827), .I2(n4826), .O(n3246) );
  AOI22S U5976 ( .A1(n4836), .A2(gray_wgt_reg[0]), .B1(n4799), .B2(
        gray_max_temp[0]), .O(n4829) );
  AOI22S U5977 ( .A1(gray_avg_reg[0]), .A2(n4854), .B1(
        SRAM_192X32_data_in_reg[24]), .B2(n4849), .O(n4828) );
  ND2S U5978 ( .I1(n4829), .I2(n4828), .O(n3243) );
  AOI22S U5979 ( .A1(n4854), .A2(gray_avg_reg[12]), .B1(n4799), .B2(
        gray_max_temp[12]), .O(n4831) );
  AOI22S U5980 ( .A1(gray_wgt_reg[12]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[20]), .B2(n4849), .O(n4830) );
  ND2S U5981 ( .I1(n4831), .I2(n4830), .O(n3247) );
  AOI22S U5982 ( .A1(n4854), .A2(gray_avg_reg[10]), .B1(n4799), .B2(
        gray_max_temp[10]), .O(n4833) );
  AOI22S U5983 ( .A1(gray_wgt_reg[10]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[18]), .B2(n4849), .O(n4832) );
  ND2S U5984 ( .I1(n4833), .I2(n4832), .O(n3249) );
  AOI22S U5985 ( .A1(n4854), .A2(gray_avg_reg[11]), .B1(n4799), .B2(
        gray_max_temp[11]), .O(n4835) );
  AOI22S U5986 ( .A1(gray_wgt_reg[11]), .A2(n4836), .B1(
        SRAM_192X32_data_in_reg[19]), .B2(n4849), .O(n4834) );
  ND2S U5987 ( .I1(n4835), .I2(n4834), .O(n3248) );
  AOI22S U5988 ( .A1(n4836), .A2(gray_wgt_reg[2]), .B1(n4854), .B2(
        gray_avg_reg[2]), .O(n4838) );
  AOI22S U5989 ( .A1(gray_max_temp[2]), .A2(n4786), .B1(
        SRAM_192X32_data_in_reg[26]), .B2(n4849), .O(n4837) );
  ND2S U5990 ( .I1(n4838), .I2(n4837), .O(n3241) );
  AOI22S U5991 ( .A1(gray_max_temp[18]), .A2(n4799), .B1(
        SRAM_192X32_data_in_reg[10]), .B2(n4849), .O(n4840) );
  AOI22S U5992 ( .A1(n4836), .A2(gray_wgt_reg[18]), .B1(n4854), .B2(
        gray_avg_reg[18]), .O(n4839) );
  ND2S U5993 ( .I1(n4840), .I2(n4839), .O(n3257) );
  AOI22S U5994 ( .A1(n4836), .A2(gray_wgt_reg[23]), .B1(n4854), .B2(
        gray_avg_reg[23]), .O(n4842) );
  AOI22S U5995 ( .A1(gray_max_temp[23]), .A2(n4786), .B1(
        SRAM_192X32_data_in_reg[15]), .B2(n4849), .O(n4841) );
  ND2S U5996 ( .I1(n4842), .I2(n4841), .O(n3252) );
  AOI22S U5997 ( .A1(gray_avg_reg[21]), .A2(n4854), .B1(
        SRAM_192X32_data_in_reg[13]), .B2(n4849), .O(n4844) );
  AOI22S U5998 ( .A1(n4836), .A2(gray_wgt_reg[21]), .B1(n4799), .B2(
        gray_max_temp[21]), .O(n4843) );
  ND2S U5999 ( .I1(n4844), .I2(n4843), .O(n3254) );
  AOI22S U6000 ( .A1(gray_max_temp[20]), .A2(n4799), .B1(
        SRAM_192X32_data_in_reg[12]), .B2(n4849), .O(n4846) );
  AOI22S U6001 ( .A1(n4836), .A2(gray_wgt_reg[20]), .B1(n4854), .B2(
        gray_avg_reg[20]), .O(n4845) );
  ND2S U6002 ( .I1(n4846), .I2(n4845), .O(n3255) );
  AOI22S U6003 ( .A1(gray_max_temp[3]), .A2(n4786), .B1(
        SRAM_192X32_data_in_reg[27]), .B2(n4849), .O(n4848) );
  AOI22S U6004 ( .A1(n4836), .A2(gray_wgt_reg[3]), .B1(n4854), .B2(
        gray_avg_reg[3]), .O(n4847) );
  ND2S U6005 ( .I1(n4848), .I2(n4847), .O(n3240) );
  AOI22S U6006 ( .A1(gray_max_temp[16]), .A2(n4799), .B1(
        SRAM_192X32_data_in_reg[8]), .B2(n4849), .O(n4851) );
  AOI22S U6007 ( .A1(n4836), .A2(gray_wgt_reg[16]), .B1(n4854), .B2(
        gray_avg_reg[16]), .O(n4850) );
  ND2S U6008 ( .I1(n4851), .I2(n4850), .O(n3259) );
  AOI22S U6009 ( .A1(gray_max_temp[7]), .A2(n4786), .B1(
        SRAM_192X32_data_in_reg[31]), .B2(n4849), .O(n4853) );
  AOI22S U6010 ( .A1(n4836), .A2(gray_wgt_reg[7]), .B1(n4854), .B2(
        gray_avg_reg[7]), .O(n4852) );
  ND2S U6011 ( .I1(n4853), .I2(n4852), .O(n3236) );
  AOI22S U6012 ( .A1(gray_max_temp[8]), .A2(n4786), .B1(
        SRAM_192X32_data_in_reg[16]), .B2(n4849), .O(n4856) );
  AOI22S U6013 ( .A1(n4836), .A2(gray_wgt_reg[8]), .B1(n4854), .B2(
        gray_avg_reg[8]), .O(n4855) );
  ND2S U6014 ( .I1(n4856), .I2(n4855), .O(n3251) );
  NR2 U6015 ( .I1(n4938), .I2(n5898), .O(n5892) );
  AOI22S U6016 ( .A1(median_in[35]), .A2(n5939), .B1(n5892), .B2(n3517), .O(
        n4860) );
  AOI22S U6017 ( .A1(median_in[43]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[91]), .O(n4859) );
  NR2 U6018 ( .I1(n4938), .I2(n4861), .O(n5901) );
  AOI22S U6019 ( .A1(median_in[36]), .A2(n5939), .B1(n5901), .B2(n3517), .O(
        n4863) );
  AOI22S U6020 ( .A1(median_in[44]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[92]), .O(n4862) );
  NR2 U6021 ( .I1(n4938), .I2(n5889), .O(n4941) );
  AOI22S U6022 ( .A1(median_in[33]), .A2(n5939), .B1(n4941), .B2(n3517), .O(
        n4865) );
  AOI22S U6023 ( .A1(median_in[41]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[89]), .O(n4864) );
  INV1S U6024 ( .I(SRAM_out_buffer[63]), .O(n6061) );
  NR2 U6025 ( .I1(n4938), .I2(n6061), .O(n5938) );
  AOI22S U6026 ( .A1(median_in[39]), .A2(n5939), .B1(n5938), .B2(n3517), .O(
        n4867) );
  AOI22S U6027 ( .A1(median_in[47]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[95]), .O(n4866) );
  INV1S U6028 ( .I(avg_temp[3]), .O(n6289) );
  NR2 U6029 ( .I1(n4871), .I2(n6289), .O(n4868) );
  MOAI1S U6030 ( .A1(n4869), .A2(n4868), .B1(n4869), .B2(avg_temp[3]), .O(
        n6204) );
  INV1S U6031 ( .I(avg_temp[2]), .O(n6293) );
  MOAI1S U6032 ( .A1(n4871), .A2(n4870), .B1(n4871), .B2(avg_temp[3]), .O(
        n6203) );
  AN2S U6033 ( .I1(n6203), .I2(avg_temp[2]), .O(n4872) );
  MOAI1S U6034 ( .A1(n6203), .A2(avg_temp[2]), .B1(n6204), .B2(n4872), .O(
        n6207) );
  MOAI1S U6035 ( .A1(n4873), .A2(n6207), .B1(n6207), .B2(avg_temp[1]), .O(
        n4874) );
  AOI22S U6036 ( .A1(median_in[54]), .A2(n6064), .B1(n4889), .B2(
        window_0__3__6_), .O(n4878) );
  AOI22S U6037 ( .A1(SRAM_out_buffer[94]), .A2(n5771), .B1(SRAM_out_buffer[86]), .B2(n4935), .O(n4877) );
  AOI22S U6038 ( .A1(median_in[55]), .A2(n6064), .B1(n4889), .B2(
        window_0__3__7_), .O(n4880) );
  AOI22S U6039 ( .A1(SRAM_out_buffer[95]), .A2(n5771), .B1(SRAM_out_buffer[87]), .B2(n4935), .O(n4879) );
  AOI22S U6040 ( .A1(window_0__4__6_), .A2(n4889), .B1(window_0__3__6_), .B2(
        n6064), .O(n4882) );
  AOI22S U6041 ( .A1(SRAM_out_buffer[86]), .A2(n5771), .B1(SRAM_out_buffer[78]), .B2(n4935), .O(n4881) );
  AOI22S U6042 ( .A1(window_0__4__7_), .A2(n4889), .B1(window_0__3__7_), .B2(
        n6064), .O(n4884) );
  AOI22S U6043 ( .A1(SRAM_out_buffer[87]), .A2(n5771), .B1(SRAM_out_buffer[79]), .B2(n4935), .O(n4883) );
  AOI22S U6044 ( .A1(window_0__4__3_), .A2(n4889), .B1(window_0__3__3_), .B2(
        n6064), .O(n4886) );
  AOI22S U6045 ( .A1(SRAM_out_buffer[83]), .A2(n5771), .B1(SRAM_out_buffer[75]), .B2(n4935), .O(n4885) );
  AOI22S U6046 ( .A1(window_0__4__1_), .A2(n4889), .B1(window_0__3__1_), .B2(
        n6064), .O(n4888) );
  AOI22S U6047 ( .A1(SRAM_out_buffer[81]), .A2(n5771), .B1(SRAM_out_buffer[73]), .B2(n4935), .O(n4887) );
  AOI22S U6048 ( .A1(window_0__4__2_), .A2(n4889), .B1(window_0__3__2_), .B2(
        n6064), .O(n4891) );
  AOI22S U6049 ( .A1(SRAM_out_buffer[82]), .A2(n5771), .B1(SRAM_out_buffer[74]), .B2(n4935), .O(n4890) );
  INV1S U6050 ( .I(SRAM_out_buffer[27]), .O(n5897) );
  INV1S U6051 ( .I(n5956), .O(n6041) );
  AOI22S U6052 ( .A1(median_in[11]), .A2(n6064), .B1(median_in[3]), .B2(n4981), 
        .O(n4895) );
  AOI22S U6053 ( .A1(median_in[51]), .A2(n6064), .B1(n4889), .B2(
        window_0__3__3_), .O(n4897) );
  AOI22S U6054 ( .A1(SRAM_out_buffer[91]), .A2(n5771), .B1(SRAM_out_buffer[83]), .B2(n4935), .O(n4896) );
  AOI22S U6055 ( .A1(median_in[52]), .A2(n6064), .B1(n4889), .B2(
        window_0__3__4_), .O(n4899) );
  AOI22S U6056 ( .A1(SRAM_out_buffer[92]), .A2(n5771), .B1(SRAM_out_buffer[84]), .B2(n4935), .O(n4898) );
  AOI22S U6057 ( .A1(median_in[49]), .A2(n6064), .B1(n4889), .B2(
        window_0__3__1_), .O(n4901) );
  AOI22S U6058 ( .A1(SRAM_out_buffer[89]), .A2(n5771), .B1(SRAM_out_buffer[81]), .B2(n4935), .O(n4900) );
  AOI22S U6059 ( .A1(median_in[53]), .A2(n6064), .B1(n4889), .B2(
        window_0__3__5_), .O(n4903) );
  AOI22S U6060 ( .A1(SRAM_out_buffer[93]), .A2(n5771), .B1(SRAM_out_buffer[85]), .B2(n4935), .O(n4902) );
  AOI22S U6061 ( .A1(window_0__4__5_), .A2(n4889), .B1(window_0__3__5_), .B2(
        n6064), .O(n4905) );
  AOI22S U6062 ( .A1(SRAM_out_buffer[85]), .A2(n5771), .B1(SRAM_out_buffer[77]), .B2(n4935), .O(n4904) );
  AOI22S U6063 ( .A1(window_0__4__0_), .A2(n4889), .B1(window_0__3__0_), .B2(
        n6064), .O(n4907) );
  AOI22S U6064 ( .A1(SRAM_out_buffer[80]), .A2(n5771), .B1(SRAM_out_buffer[72]), .B2(n4935), .O(n4906) );
  AOI22S U6065 ( .A1(window_0__4__4_), .A2(n4889), .B1(window_0__3__4_), .B2(
        n6064), .O(n4909) );
  AOI22S U6066 ( .A1(SRAM_out_buffer[84]), .A2(n5771), .B1(SRAM_out_buffer[76]), .B2(n4935), .O(n4908) );
  AOI22S U6067 ( .A1(median_in[38]), .A2(n5939), .B1(n5925), .B2(n3517), .O(
        n4911) );
  AOI22S U6068 ( .A1(median_in[46]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[94]), .O(n4910) );
  AOI22S U6069 ( .A1(median_in[37]), .A2(n5939), .B1(n5912), .B2(n3517), .O(
        n4913) );
  AOI22S U6070 ( .A1(median_in[45]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[93]), .O(n4912) );
  AOI22S U6071 ( .A1(median_in[32]), .A2(n5939), .B1(n4917), .B2(n3517), .O(
        n4916) );
  AOI22S U6072 ( .A1(median_in[40]), .A2(n6064), .B1(n4971), .B2(
        SRAM_out_buffer[88]), .O(n4915) );
  INV1S U6073 ( .I(median_in[32]), .O(n5207) );
  MOAI1S U6074 ( .A1(n5942), .A2(n5207), .B1(SRAM_out_buffer[88]), .B2(n5935), 
        .O(n4919) );
  NR2 U6075 ( .I1(n5176), .I2(n5943), .O(n4918) );
  INV1S U6076 ( .I(n6114), .O(n4920) );
  FA1 U6077 ( .A(N1046), .B(n4923), .CI(n4922), .CO(n5114), .S(n4738) );
  ND2S U6078 ( .I1(n4924), .I2(n5131), .O(n4927) );
  AOI22S U6079 ( .A1(n5126), .A2(SRAM_64X32_addr[4]), .B1(n5124), .B2(N1047), 
        .O(n4926) );
  ND3S U6080 ( .I1(n4927), .I2(n4926), .I3(n4925), .O(n2592) );
  INV1S U6081 ( .I(n4935), .O(n5941) );
  INV1S U6082 ( .I(SRAM_out_buffer[90]), .O(n4933) );
  INV1S U6083 ( .I(median_in[50]), .O(n5528) );
  OAI222S U6084 ( .A1(n5941), .A2(n4933), .B1(n5527), .B2(n5942), .C1(n5528), 
        .C2(n5943), .O(n2980) );
  ND2S U6085 ( .I1(n5725), .I2(n6243), .O(n4930) );
  AO13S U6086 ( .B1(n4932), .B2(n4931), .B3(n4930), .A1(n4929), .O(n5946) );
  OAI222S U6087 ( .A1(n5943), .A2(n5527), .B1(n5533), .B2(n5942), .C1(n4933), 
        .C2(n5946), .O(n2979) );
  INV1S U6088 ( .I(SRAM_out_buffer[88]), .O(n4934) );
  OAI222S U6089 ( .A1(n5943), .A2(n5524), .B1(n5545), .B2(n5942), .C1(n4934), 
        .C2(n5946), .O(n3003) );
  INV1S U6090 ( .I(SRAM_out_buffer[89]), .O(n4936) );
  OAI222S U6091 ( .A1(n5943), .A2(n5525), .B1(n5534), .B2(n5942), .C1(n4936), 
        .C2(n5946), .O(n2991) );
  NR2 U6092 ( .I1(n4938), .I2(n4937), .O(n4970) );
  MOAI1S U6093 ( .A1(n5942), .A2(n5178), .B1(n5935), .B2(SRAM_out_buffer[90]), 
        .O(n4939) );
  MOAI1S U6094 ( .A1(n5942), .A2(n5177), .B1(n5935), .B2(SRAM_out_buffer[89]), 
        .O(n4940) );
  NR2 U6095 ( .I1(n4942), .I2(n5709), .O(n4944) );
  NR2 U6096 ( .I1(n5695), .I2(n4944), .O(n4946) );
  NR2 U6097 ( .I1(n4969), .I2(n4943), .O(n4966) );
  MOAI1S U6098 ( .A1(n4946), .A2(n4945), .B1(n4944), .B2(n4966), .O(n3223) );
  NR2 U6099 ( .I1(n4947), .I2(n3517), .O(n4962) );
  INV1S U6100 ( .I(conv_dly3[2]), .O(n5594) );
  ND3S U6101 ( .I1(conv_dly3[0]), .I2(conv_dly3[1]), .I3(n5594), .O(n5593) );
  ND2S U6102 ( .I1(n4956), .I2(n5593), .O(n4955) );
  OA12S U6103 ( .B1(n4952), .B2(n4948), .A1(n4955), .O(n4953) );
  INV1S U6104 ( .I(n4952), .O(n4958) );
  AOI13HS U6105 ( .B1(n4958), .B2(n6069), .B3(N6291), .A1(
        wait_conv_out_count[3]), .O(n4950) );
  INV1S U6106 ( .I(n5593), .O(n4949) );
  ND2S U6107 ( .I1(n5591), .I2(n4949), .O(n4959) );
  OAI12HS U6108 ( .B1(n4953), .B2(n4950), .A1(n4959), .O(n3363) );
  OAI22S U6109 ( .A1(n5105), .A2(n4953), .B1(n4952), .B2(n4951), .O(n3366) );
  ND2S U6110 ( .I1(n4958), .I2(n6302), .O(n4954) );
  OAI112HS U6111 ( .C1(n6302), .C2(n4955), .A1(n4954), .B1(n5591), .O(n3365)
         );
  INV1S U6112 ( .I(n4956), .O(n5596) );
  ND3S U6113 ( .I1(n4958), .I2(n4957), .I3(n6071), .O(n4960) );
  OAI112HS U6114 ( .C1(n5596), .C2(n6070), .A1(n4960), .B1(n4959), .O(n3367)
         );
  ND2S U6115 ( .I1(n5596), .I2(n6069), .O(n4965) );
  ND2S U6116 ( .I1(n4962), .I2(n4961), .O(n4963) );
  ND3S U6117 ( .I1(n4963), .I2(n5593), .I3(n5591), .O(n4964) );
  AO12S U6118 ( .B1(n4965), .B2(N6291), .A1(n4964), .O(n3364) );
  NR2 U6119 ( .I1(n4966), .I2(n5709), .O(n4968) );
  MOAI1S U6120 ( .A1(n6301), .A2(n4969), .B1(n4968), .B2(n4967), .O(n3222) );
  INV1S U6121 ( .I(n5709), .O(n5715) );
  AOI22S U6122 ( .A1(n6064), .A2(median_in[42]), .B1(n4971), .B2(
        SRAM_out_buffer[90]), .O(n4972) );
  OAI112HS U6123 ( .C1(n5943), .C2(n5178), .A1(n4973), .B1(n4972), .O(n2982)
         );
  ND2S U6124 ( .I1(median_in[17]), .I2(n6064), .O(n4974) );
  AOI22S U6125 ( .A1(median_in[11]), .A2(n4981), .B1(n6064), .B2(median_in[19]), .O(n4979) );
  OAI12HS U6126 ( .B1(n4980), .B2(n5918), .A1(n4979), .O(n2963) );
  AOI22S U6127 ( .A1(median_in[16]), .A2(n6064), .B1(median_in[8]), .B2(n4981), 
        .O(n4982) );
  OAI112HS U6128 ( .C1(n4984), .C2(n5918), .A1(n4983), .B1(n4982), .O(n2999)
         );
  INV1S U6129 ( .I(SRAM_out_buffer[92]), .O(n5903) );
  OAI222S U6130 ( .A1(n5532), .A2(n5942), .B1(n5943), .B2(n5902), .C1(n5903), 
        .C2(n5946), .O(n2955) );
  NR2 U6131 ( .I1(n6015), .I2(n4985), .O(n4987) );
  OA12S U6132 ( .B1(cal_count_5[0]), .B2(n6301), .A1(n5711), .O(n3215) );
  INV1S U6133 ( .I(in_valid2), .O(n5572) );
  MOAI1S U6134 ( .A1(n5009), .A2(n3533), .B1(n4991), .B2(n5006), .O(n2604) );
  INV1S U6135 ( .I(N1047), .O(n4994) );
  MOAI1S U6136 ( .A1(n4994), .A2(n5009), .B1(n4993), .B2(n5006), .O(n2602) );
  INV1S U6137 ( .I(N1046), .O(n4997) );
  MOAI1S U6138 ( .A1(n4997), .A2(n5009), .B1(n4996), .B2(n5006), .O(n2601) );
  INV1S U6139 ( .I(N1045), .O(n5001) );
  MOAI1S U6140 ( .A1(n5009), .A2(n5001), .B1(n5000), .B2(n5006), .O(n2600) );
  INV1S U6141 ( .I(rd_addr[7]), .O(n5008) );
  XOR2HS U6142 ( .I1(rd_addr[7]), .I2(n5003), .O(n5005) );
  FA1S U6143 ( .A(rd_addr[6]), .B(n5003), .CI(n5002), .CO(n5004), .S(n4991) );
  XOR2HS U6144 ( .I1(n5005), .I2(n5004), .O(n5007) );
  MOAI1S U6145 ( .A1(n5009), .A2(n5008), .B1(n5007), .B2(n5006), .O(n2605) );
  INV1S U6146 ( .I(wb_addr[2]), .O(n5054) );
  ND2S U6147 ( .I1(wb_addr[0]), .I2(wb_addr[1]), .O(n5051) );
  NR2 U6148 ( .I1(n5054), .I2(n5051), .O(n5050) );
  ND2S U6149 ( .I1(wb_addr[3]), .I2(n5050), .O(n5038) );
  NR2 U6150 ( .I1(n5041), .I2(n5038), .O(n5037) );
  ND2S U6151 ( .I1(wb_addr[5]), .I2(n5037), .O(n5017) );
  AN2B1S U6152 ( .I1(wb_addr[6]), .B1(n5017), .O(n5012) );
  AOI13HS U6153 ( .B1(n5582), .B2(n3647), .B3(n6245), .A1(n6300), .O(n5011) );
  INV1S U6154 ( .I(n5055), .O(n5064) );
  NR2 U6155 ( .I1(n5013), .I2(n5064), .O(n5063) );
  OAI12HS U6156 ( .B1(n5013), .B2(n5012), .A1(n5055), .O(n5016) );
  INV1S U6157 ( .I(n5063), .O(n5066) );
  OAI12HS U6158 ( .B1(wb_addr[5]), .B2(n5037), .A1(n5017), .O(n5015) );
  MOAI1S U6159 ( .A1(n5066), .A2(n5015), .B1(wb_addr[5]), .B2(n5064), .O(n3199) );
  ND2S U6160 ( .I1(n5063), .I2(n5016), .O(n5018) );
  MOAI1S U6161 ( .A1(n5018), .A2(n5017), .B1(n5016), .B2(wb_addr[6]), .O(n3198) );
  XNR2HS U6162 ( .I1(n5020), .I2(n5019), .O(n5022) );
  XNR2HS U6163 ( .I1(n5022), .I2(n5021), .O(n5023) );
  ND2S U6164 ( .I1(n5023), .I2(n5098), .O(n5029) );
  OA112S U6165 ( .C1(n5098), .C2(n6303), .A1(n5025), .B1(n5095), .O(n5028) );
  ND3S U6166 ( .I1(n5029), .I2(n5028), .I3(n5027), .O(n3206) );
  ND3S U6167 ( .I1(n5034), .I2(n5095), .I3(n5033), .O(n5035) );
  NR2 U6168 ( .I1(n5037), .I2(n5066), .O(n5040) );
  ND2S U6169 ( .I1(n5041), .I2(n5038), .O(n5039) );
  MOAI1S U6170 ( .A1(n5055), .A2(n5041), .B1(n5040), .B2(n5039), .O(n3200) );
  XNR2HS U6171 ( .I1(n5050), .I2(wb_addr[3]), .O(n5042) );
  MOAI1S U6172 ( .A1(n5066), .A2(n5042), .B1(wb_addr[3]), .B2(n5064), .O(n3201) );
  FA1 U6173 ( .A(n5045), .B(n5044), .CI(n5043), .CO(n5089), .S(n5049) );
  ND3S U6174 ( .I1(n5047), .I2(n5095), .I3(n5046), .O(n5048) );
  NR2 U6175 ( .I1(n5050), .I2(n5066), .O(n5053) );
  ND2S U6176 ( .I1(n5054), .I2(n5051), .O(n5052) );
  MOAI1S U6177 ( .A1(n5055), .A2(n5054), .B1(n5053), .B2(n5052), .O(n3202) );
  FA1 U6178 ( .A(n5058), .B(n5057), .CI(n5056), .CO(n5043), .S(n5062) );
  ND3S U6179 ( .I1(n5060), .I2(n5095), .I3(n5059), .O(n5061) );
  XNR2HS U6180 ( .I1(wb_addr[0]), .I2(wb_addr[1]), .O(n5065) );
  MOAI1S U6181 ( .A1(n5066), .A2(n5065), .B1(wb_addr[1]), .B2(n5064), .O(n3203) );
  ND2S U6182 ( .I1(n5068), .I2(n5067), .O(n5077) );
  FA1 U6183 ( .A(n5071), .B(n5070), .CI(n5069), .CO(n5056), .S(n5072) );
  OR2S U6184 ( .I1(n3506), .I2(n5072), .O(n5076) );
  ND3S U6185 ( .I1(n5074), .I2(n5095), .I3(n5073), .O(n5075) );
  NR2 U6186 ( .I1(n3486), .I2(n5077), .O(n5078) );
  XOR2HS U6187 ( .I1(n5080), .I2(n5079), .O(n5081) );
  XNR2HS U6188 ( .I1(n5082), .I2(n5081), .O(n5083) );
  OR2S U6189 ( .I1(n5084), .I2(n5083), .O(n5088) );
  ND3S U6190 ( .I1(n5086), .I2(n5095), .I3(n5085), .O(n5087) );
  FA1 U6191 ( .A(n5091), .B(n5090), .CI(n5089), .CO(n5030), .S(n5099) );
  ND3S U6192 ( .I1(n5096), .I2(n5095), .I3(n5094), .O(n5097) );
  INV1S U6193 ( .I(template_count[2]), .O(n5102) );
  NR2 U6194 ( .I1(n5102), .I2(n5100), .O(n5631) );
  INV1S U6195 ( .I(n5100), .O(n5629) );
  NR2 U6196 ( .I1(template_count[0]), .I2(template_count[1]), .O(n5103) );
  INV1S U6197 ( .I(template_count[0]), .O(n5632) );
  NR2 U6198 ( .I1(template_count[1]), .I2(n5632), .O(n5636) );
  INV1S U6199 ( .I(n5633), .O(n5635) );
  AOI13HS U6200 ( .B1(n5106), .B2(n61150), .B3(n5105), .A1(out_valid), .O(
        n61190) );
  NR2 U6201 ( .I1(n61190), .I2(n61230), .O(n3196) );
  FA1 U6202 ( .A(N1044), .B(n5108), .CI(n5107), .CO(n4736), .S(n5113) );
  ND2S U6203 ( .I1(SRAM_64X32_addr[1]), .I2(n5126), .O(n5111) );
  AOI22S U6204 ( .A1(N1044), .A2(n5124), .B1(wb_addr[1]), .B2(n5123), .O(n5110) );
  XOR2HS U6205 ( .I1(N1048), .I2(n5122), .O(n5116) );
  FA1 U6206 ( .A(N1047), .B(n5122), .CI(n5114), .CO(n5115), .S(n4924) );
  XOR2HS U6207 ( .I1(n5116), .I2(n5115), .O(n5117) );
  ND2S U6208 ( .I1(n5117), .I2(n5131), .O(n5120) );
  AOI22S U6209 ( .A1(n5126), .A2(SRAM_64X32_addr[5]), .B1(n5124), .B2(N1048), 
        .O(n5119) );
  ND3S U6210 ( .I1(n5120), .I2(n5119), .I3(n5118), .O(n2591) );
  FA1 U6211 ( .A(n5122), .B(N1043), .CI(n5121), .CO(n5107), .S(n5132) );
  OAI22S U6212 ( .A1(n5126), .A2(n5125), .B1(SRAM_64X32_addr[0]), .B2(n5125), 
        .O(n5127) );
  NR2 U6213 ( .I1(n5135), .I2(n5610), .O(N813) );
  NR2 U6214 ( .I1(n5135), .I2(n5134), .O(N814) );
  FA1S U6215 ( .A(median_in[25]), .B(median_in[24]), .CI(n5177), .CO(n5136) );
  FA1S U6216 ( .A(n5178), .B(median_in[26]), .CI(n5136), .CO(n5137) );
  FA1S U6217 ( .A(n5890), .B(median_in[27]), .CI(n5137), .CO(n5138) );
  FA1S U6218 ( .A(n5899), .B(median_in[28]), .CI(n5138), .CO(n5139) );
  ND2S U6219 ( .I1(median_in[35]), .I2(n5186), .O(n5147) );
  OAI12HS U6220 ( .B1(n5144), .B2(n5143), .A1(n5142), .O(n5146) );
  AOI13HS U6221 ( .B1(n5148), .B2(n5147), .B3(n5146), .A1(n5145), .O(n5150) );
  OAI22S U6222 ( .A1(n5150), .A2(n5149), .B1(n5205), .B2(median_in[39]), .O(
        n5160) );
  MOAI1 U6223 ( .A1(n5151), .A2(n5187), .B1(n5151), .B2(n5160), .O(n5180) );
  MOAI1S U6224 ( .A1(n5183), .A2(median_in[30]), .B1(median_in[47]), .B2(n5206), .O(n5168) );
  INV1S U6225 ( .I(n5168), .O(n5161) );
  AOI22S U6226 ( .A1(median_in[26]), .A2(n6313), .B1(median_in[27]), .B2(n5186), .O(n5163) );
  INV1S U6227 ( .I(median_in[41]), .O(n5188) );
  MOAI1S U6228 ( .A1(n5188), .A2(median_in[25]), .B1(median_in[42]), .B2(n6318), .O(n5165) );
  OR2S U6229 ( .I1(n5165), .I2(median_in[40]), .O(n5155) );
  ND2S U6230 ( .I1(median_in[42]), .I2(n6318), .O(n5152) );
  ND3S U6231 ( .I1(median_in[25]), .I2(n5188), .I3(n5152), .O(n5154) );
  AOI22S U6232 ( .A1(median_in[43]), .A2(n6319), .B1(median_in[44]), .B2(n6311), .O(n5153) );
  ND2S U6233 ( .I1(median_in[45]), .I2(n5179), .O(n5158) );
  ND2S U6234 ( .I1(n5153), .I2(n5158), .O(n5167) );
  AOI13HS U6235 ( .B1(n5163), .B2(n5155), .B3(n5154), .A1(n5167), .O(n5156) );
  NR2 U6236 ( .I1(n5156), .I2(n5160), .O(n5159) );
  MOAI1S U6237 ( .A1(n5179), .A2(median_in[45]), .B1(n5183), .B2(median_in[30]), .O(n5157) );
  AOI13HS U6238 ( .B1(median_in[28]), .B2(n5185), .B3(n5158), .A1(n5157), .O(
        n5170) );
  MOAI1S U6239 ( .A1(n5161), .A2(n5160), .B1(n5159), .B2(n5170), .O(n5174) );
  NR2 U6240 ( .I1(median_in[41]), .I2(n6310), .O(n5162) );
  NR2 U6241 ( .I1(median_in[24]), .I2(n5162), .O(n5164) );
  OAI12HS U6242 ( .B1(n5165), .B2(n5164), .A1(n5163), .O(n5166) );
  OR2B1S U6243 ( .I1(n5167), .B1(n5166), .O(n5169) );
  AOI22S U6244 ( .A1(n5174), .A2(n5173), .B1(n5172), .B2(n5187), .O(n5181) );
  OAI222S U6245 ( .A1(n5182), .A2(n5176), .B1(n5207), .B2(n5180), .C1(n5175), 
        .C2(n5181), .O(find_median_inst_mid2[0]) );
  OAI222S U6246 ( .A1(n5182), .A2(n6310), .B1(n5188), .B2(n5181), .C1(n5177), 
        .C2(n5180), .O(find_median_inst_mid2[1]) );
  OAI222S U6247 ( .A1(n5182), .A2(n6318), .B1(n6313), .B2(n5181), .C1(n5178), 
        .C2(n5180), .O(find_median_inst_mid2[2]) );
  OAI222S U6248 ( .A1(n5182), .A2(n6319), .B1(n5186), .B2(n5181), .C1(n5890), 
        .C2(n5180), .O(find_median_inst_mid2[3]) );
  OAI222S U6249 ( .A1(n5182), .A2(n6311), .B1(n5185), .B2(n5181), .C1(n5899), 
        .C2(n5180), .O(find_median_inst_mid2[4]) );
  OAI222S U6250 ( .A1(n5182), .A2(n5179), .B1(n5184), .B2(n5181), .C1(n5910), 
        .C2(n5180), .O(find_median_inst_mid2[5]) );
  OAI222S U6251 ( .A1(n5182), .A2(n6312), .B1(n5923), .B2(n5180), .C1(n5183), 
        .C2(n5181), .O(find_median_inst_mid2[6]) );
  OAI222S U6252 ( .A1(n5182), .A2(n5206), .B1(n5205), .B2(n5181), .C1(n5936), 
        .C2(n5180), .O(find_median_inst_mid2[7]) );
  MOAI1S U6253 ( .A1(n5208), .A2(median_in[38]), .B1(n5208), .B2(n5183), .O(
        n5203) );
  MOAI1S U6254 ( .A1(n5208), .A2(median_in[37]), .B1(n5208), .B2(n5184), .O(
        n5202) );
  MOAI1S U6255 ( .A1(n5208), .A2(median_in[36]), .B1(n5208), .B2(n5185), .O(
        n5201) );
  MOAI1S U6256 ( .A1(n5208), .A2(median_in[35]), .B1(n5208), .B2(n5186), .O(
        n5200) );
  MOAI1S U6257 ( .A1(n5208), .A2(median_in[34]), .B1(n5208), .B2(n6313), .O(
        n5199) );
  MOAI1S U6258 ( .A1(n5187), .A2(median_in[40]), .B1(n5187), .B2(n5207), .O(
        n5197) );
  FA1S U6259 ( .A(n5197), .B(median_in[25]), .CI(n5198), .CO(n5189) );
  FA1S U6260 ( .A(median_in[26]), .B(n5199), .CI(n5189), .CO(n5190) );
  FA1S U6261 ( .A(n5200), .B(median_in[27]), .CI(n5190), .CO(n5191) );
  FA1S U6262 ( .A(median_in[28]), .B(n5201), .CI(n5191), .CO(n5192) );
  FA1S U6263 ( .A(n5202), .B(median_in[29]), .CI(n5192), .CO(n5193) );
  MOAI1S U6264 ( .A1(n5204), .A2(n5197), .B1(n5204), .B2(median_in[24]), .O(
        find_median_inst_min2[0]) );
  MOAI1S U6265 ( .A1(n5204), .A2(n5198), .B1(n5204), .B2(median_in[25]), .O(
        find_median_inst_min2[1]) );
  MOAI1S U6266 ( .A1(n5204), .A2(n5199), .B1(n5204), .B2(median_in[26]), .O(
        find_median_inst_min2[2]) );
  MOAI1S U6267 ( .A1(n5204), .A2(n5200), .B1(n5204), .B2(median_in[27]), .O(
        find_median_inst_min2[3]) );
  MOAI1S U6268 ( .A1(n5204), .A2(n5201), .B1(n5204), .B2(median_in[28]), .O(
        find_median_inst_min2[4]) );
  MOAI1S U6269 ( .A1(n5204), .A2(n5202), .B1(n5204), .B2(median_in[29]), .O(
        find_median_inst_min2[5]) );
  MOAI1S U6270 ( .A1(n5204), .A2(n5203), .B1(n5204), .B2(median_in[30]), .O(
        find_median_inst_min2[6]) );
  NR3 U6271 ( .I1(n5936), .I2(n5206), .I3(n5205), .O(find_median_inst_min2[7])
         );
  MOAI1S U6272 ( .A1(n5208), .A2(median_in[40]), .B1(n5208), .B2(n5207), .O(
        n5209) );
  MOAI1S U6273 ( .A1(n5211), .A2(n5209), .B1(n5211), .B2(median_in[24]), .O(
        find_median_inst_max2[0]) );
  MOAI1S U6274 ( .A1(n5211), .A2(n5210), .B1(n5211), .B2(median_in[29]), .O(
        find_median_inst_max2[5]) );
  ND2S U6275 ( .I1(median_in[5]), .I2(n5922), .O(n5218) );
  ND2S U6276 ( .I1(median_in[13]), .I2(n5269), .O(n5215) );
  NR2 U6277 ( .I1(n5221), .I2(n5220), .O(n5222) );
  NR2 U6278 ( .I1(median_in[17]), .I2(n5263), .O(n5224) );
  NR2 U6279 ( .I1(n5224), .I2(n5226), .O(n5225) );
  INV1S U6280 ( .I(median_in[8]), .O(n5261) );
  MOAI1S U6281 ( .A1(n5227), .A2(n5226), .B1(n5225), .B2(n5261), .O(n5230) );
  OAI12HS U6282 ( .B1(n5230), .B2(n5229), .A1(n5228), .O(n5231) );
  MOAI1S U6283 ( .A1(n6067), .A2(median_in[23]), .B1(n5232), .B2(n5231), .O(
        n5257) );
  MOAI1 U6284 ( .A1(n5234), .A2(n5257), .B1(n5234), .B2(n5233), .O(n5272) );
  ND2S U6285 ( .I1(median_in[21]), .I2(n5269), .O(n5237) );
  NR2 U6286 ( .I1(median_in[21]), .I2(n5269), .O(n5235) );
  AOI13HS U6287 ( .B1(median_in[4]), .B2(n5909), .B3(n5237), .A1(n5235), .O(
        n5251) );
  NR2 U6288 ( .I1(median_in[17]), .I2(n6314), .O(n5244) );
  AOI22S U6289 ( .A1(median_in[17]), .A2(n6314), .B1(median_in[18]), .B2(n6315), .O(n5247) );
  OA12S U6290 ( .B1(median_in[0]), .B2(n5244), .A1(n5247), .O(n5238) );
  MOAI1S U6291 ( .A1(n6316), .A2(median_in[19]), .B1(n5266), .B2(median_in[2]), 
        .O(n5245) );
  MOAI1S U6292 ( .A1(median_in[3]), .A2(n5268), .B1(n6317), .B2(median_in[20]), 
        .O(n5236) );
  AN2B1S U6293 ( .I1(n5237), .B1(n5236), .O(n5249) );
  OAI12HS U6294 ( .B1(n5238), .B2(n5245), .A1(n5249), .O(n5239) );
  AOI22S U6295 ( .A1(median_in[22]), .A2(n6322), .B1(n5251), .B2(n5239), .O(
        n5240) );
  NR2 U6296 ( .I1(n5240), .I2(n5252), .O(n5241) );
  NR2 U6297 ( .I1(n5243), .I2(n5241), .O(n5258) );
  NR2 U6298 ( .I1(median_in[6]), .I2(n5271), .O(n5242) );
  NR2 U6299 ( .I1(n5243), .I2(n5242), .O(n5254) );
  OR2S U6300 ( .I1(n5260), .I2(n5244), .O(n5246) );
  AO12S U6301 ( .B1(n5247), .B2(n5246), .A1(n5245), .O(n5248) );
  ND2S U6302 ( .I1(n5249), .I2(n5248), .O(n5250) );
  ND2S U6303 ( .I1(n5251), .I2(n5250), .O(n5253) );
  OAI22S U6304 ( .A1(n5255), .A2(n5254), .B1(n5253), .B2(n5252), .O(n5256) );
  AOI22S U6305 ( .A1(n5259), .A2(n5258), .B1(n5257), .B2(n5256), .O(n5273) );
  OAI222S U6306 ( .A1(n5274), .A2(n5262), .B1(n5261), .B2(n5272), .C1(n5260), 
        .C2(n5273), .O(find_median_inst_mid3[0]) );
  OAI222S U6307 ( .A1(n5274), .A2(n6314), .B1(n5264), .B2(n5273), .C1(n5263), 
        .C2(n5272), .O(find_median_inst_mid3[1]) );
  OAI222S U6308 ( .A1(n5274), .A2(n6315), .B1(n5266), .B2(n5273), .C1(n5265), 
        .C2(n5272), .O(find_median_inst_mid3[2]) );
  OAI222S U6309 ( .A1(n5274), .A2(n6316), .B1(n5268), .B2(n5273), .C1(n5267), 
        .C2(n5272), .O(find_median_inst_mid3[3]) );
  OAI222S U6310 ( .A1(n5274), .A2(n6317), .B1(n5909), .B2(n5273), .C1(n5906), 
        .C2(n5272), .O(find_median_inst_mid3[4]) );
  OAI222S U6311 ( .A1(n5274), .A2(n5269), .B1(n5919), .B2(n5273), .C1(n5922), 
        .C2(n5272), .O(find_median_inst_mid3[5]) );
  OAI222S U6312 ( .A1(n5274), .A2(n6322), .B1(n5271), .B2(n5273), .C1(n5270), 
        .C2(n5272), .O(find_median_inst_mid3[6]) );
  OAI222S U6313 ( .A1(n5274), .A2(n5276), .B1(n5275), .B2(n5273), .C1(n6067), 
        .C2(n5272), .O(find_median_inst_mid3[7]) );
  NR3 U6314 ( .I1(n6067), .I2(n5276), .I3(n5275), .O(find_median_inst_min3[7])
         );
  MOAI1S U6315 ( .A1(n5279), .A2(n5277), .B1(n5279), .B2(median_in[0]), .O(
        find_median_inst_max3[0]) );
  MOAI1S U6316 ( .A1(n5279), .A2(n5278), .B1(n5279), .B2(median_in[5]), .O(
        find_median_inst_max3[5]) );
  INV1S U6317 ( .I(find_median_inst_max1_reg[7]), .O(n5292) );
  INV1S U6318 ( .I(find_median_inst_max1_reg[6]), .O(n5290) );
  INV1S U6319 ( .I(find_median_inst_max1_reg[5]), .O(n5288) );
  INV1S U6320 ( .I(find_median_inst_max1_reg[4]), .O(n5286) );
  INV1S U6321 ( .I(find_median_inst_max1_reg[3]), .O(n5284) );
  INV1S U6322 ( .I(find_median_inst_max1_reg[2]), .O(n5282) );
  INV1S U6323 ( .I(find_median_inst_max1_reg[1]), .O(n5280) );
  OAI22S U6324 ( .A1(n5293), .A2(find_median_inst_max2_reg[6]), .B1(n5294), 
        .B2(find_median_inst_max1_reg[6]), .O(n5311) );
  AOI22S U6325 ( .A1(n5294), .A2(find_median_inst_max2_reg[5]), .B1(n5293), 
        .B2(find_median_inst_max1_reg[5]), .O(n5310) );
  OAI22S U6326 ( .A1(n5293), .A2(find_median_inst_max2_reg[4]), .B1(n5294), 
        .B2(find_median_inst_max1_reg[4]), .O(n5309) );
  OAI22S U6327 ( .A1(n5293), .A2(find_median_inst_max2_reg[3]), .B1(n5294), 
        .B2(find_median_inst_max1_reg[3]), .O(n5308) );
  OAI22S U6328 ( .A1(n5293), .A2(find_median_inst_max2_reg[2]), .B1(n5294), 
        .B2(find_median_inst_max1_reg[2]), .O(n5307) );
  OAI22S U6329 ( .A1(n5293), .A2(find_median_inst_max2_reg[1]), .B1(n5294), 
        .B2(find_median_inst_max1_reg[1]), .O(n5306) );
  OAI22S U6330 ( .A1(n5294), .A2(find_median_inst_max1_reg[0]), .B1(n5293), 
        .B2(find_median_inst_max2_reg[0]), .O(n5305) );
  NR2 U6331 ( .I1(n5299), .I2(n5298), .O(n5301) );
  NR2 U6332 ( .I1(find_median_inst_max3_reg[5]), .I2(n5310), .O(n5300) );
  NR2 U6333 ( .I1(n5301), .I2(n5300), .O(n5302) );
  ND2S U6334 ( .I1(find_median_inst_max3_reg[7]), .I2(n5304), .O(n5303) );
  MOAI1S U6335 ( .A1(n5312), .A2(n5305), .B1(n5312), .B2(
        find_median_inst_max3_reg[0]), .O(find_median_inst_max_min[0]) );
  MOAI1S U6336 ( .A1(n5312), .A2(n5306), .B1(n5312), .B2(
        find_median_inst_max3_reg[1]), .O(find_median_inst_max_min[1]) );
  MOAI1S U6337 ( .A1(n5312), .A2(n5307), .B1(n5312), .B2(
        find_median_inst_max3_reg[2]), .O(find_median_inst_max_min[2]) );
  MOAI1S U6338 ( .A1(n5312), .A2(n5308), .B1(n5312), .B2(
        find_median_inst_max3_reg[3]), .O(find_median_inst_max_min[3]) );
  MOAI1S U6339 ( .A1(n5312), .A2(n5309), .B1(n5312), .B2(
        find_median_inst_max3_reg[4]), .O(find_median_inst_max_min[4]) );
  MOAI1S U6340 ( .A1(n5312), .A2(n5310), .B1(n5312), .B2(
        find_median_inst_max3_reg[5]), .O(find_median_inst_max_min[5]) );
  MOAI1S U6341 ( .A1(n5312), .A2(n5311), .B1(n5312), .B2(
        find_median_inst_max3_reg[6]), .O(find_median_inst_max_min[6]) );
  AN2S U6342 ( .I1(n5313), .I2(find_median_inst_max3_reg[7]), .O(
        find_median_inst_max_min[7]) );
  INV1S U6343 ( .I(find_median_inst_mid3_reg[4]), .O(n5362) );
  INV1S U6344 ( .I(find_median_inst_mid2_reg[5]), .O(n5379) );
  NR2 U6345 ( .I1(n5379), .I2(find_median_inst_mid3_reg[5]), .O(n5314) );
  ND2S U6346 ( .I1(n5379), .I2(find_median_inst_mid3_reg[5]), .O(n5315) );
  OA13S U6347 ( .B1(n5362), .B2(find_median_inst_mid2_reg[4]), .B3(n5314), 
        .A1(n5315), .O(n5345) );
  INV1S U6348 ( .I(find_median_inst_mid2_reg[6]), .O(n5385) );
  ND2S U6349 ( .I1(find_median_inst_mid3_reg[6]), .I2(n5385), .O(n5319) );
  INV1S U6350 ( .I(find_median_inst_mid2_reg[3]), .O(n5377) );
  ND2S U6351 ( .I1(find_median_inst_mid3_reg[3]), .I2(n5377), .O(n5344) );
  INV1S U6352 ( .I(find_median_inst_mid2_reg[2]), .O(n5374) );
  ND2S U6353 ( .I1(find_median_inst_mid3_reg[2]), .I2(n5374), .O(n5341) );
  INV1S U6354 ( .I(find_median_inst_mid3_reg[1]), .O(n5358) );
  NR2 U6355 ( .I1(find_median_inst_mid2_reg[1]), .I2(n5358), .O(n5343) );
  ND2S U6356 ( .I1(find_median_inst_mid2_reg[1]), .I2(n5358), .O(n5340) );
  INV1S U6357 ( .I(find_median_inst_mid3_reg[2]), .O(n5375) );
  ND2S U6358 ( .I1(find_median_inst_mid2_reg[2]), .I2(n5375), .O(n5350) );
  OAI112HS U6359 ( .C1(find_median_inst_mid3_reg[0]), .C2(n5343), .A1(n5340), 
        .B1(n5350), .O(n5317) );
  AOI13HS U6360 ( .B1(find_median_inst_mid2_reg[4]), .B2(n5362), .B3(n5315), 
        .A1(n5314), .O(n5347) );
  OA12S U6361 ( .B1(find_median_inst_mid3_reg[3]), .B2(n5377), .A1(n5347), .O(
        n5351) );
  INV1S U6362 ( .I(n5351), .O(n5316) );
  AO13S U6363 ( .B1(n5344), .B2(n5341), .B3(n5317), .A1(n5316), .O(n5318) );
  INV1S U6364 ( .I(find_median_inst_mid2_reg[7]), .O(n5352) );
  OAI22S U6365 ( .A1(find_median_inst_mid3_reg[7]), .A2(n5352), .B1(n5385), 
        .B2(find_median_inst_mid3_reg[6]), .O(n5353) );
  AOI13HS U6366 ( .B1(n5345), .B2(n5319), .B3(n5318), .A1(n5353), .O(n5357) );
  INV1S U6367 ( .I(find_median_inst_mid1_reg[3]), .O(n5376) );
  INV1S U6368 ( .I(find_median_inst_mid1_reg[2]), .O(n5373) );
  INV1S U6369 ( .I(find_median_inst_mid1_reg[1]), .O(n5320) );
  INV1S U6370 ( .I(find_median_inst_mid1_reg[5]), .O(n5380) );
  ND2S U6371 ( .I1(n5380), .I2(find_median_inst_mid2_reg[5]), .O(n5323) );
  INV1S U6372 ( .I(find_median_inst_mid2_reg[4]), .O(n5325) );
  NR2 U6373 ( .I1(n5380), .I2(find_median_inst_mid2_reg[5]), .O(n5324) );
  AOI13HS U6374 ( .B1(find_median_inst_mid1_reg[4]), .B2(n5323), .B3(n5325), 
        .A1(n5324), .O(n5334) );
  ND2S U6375 ( .I1(n5332), .I2(n5334), .O(n5326) );
  OA13S U6376 ( .B1(n5325), .B2(n5324), .B3(find_median_inst_mid1_reg[4]), 
        .A1(n5323), .O(n5331) );
  INV1S U6377 ( .I(find_median_inst_mid1_reg[6]), .O(n5383) );
  ND2S U6378 ( .I1(find_median_inst_mid2_reg[6]), .I2(n5383), .O(n5338) );
  INV1S U6379 ( .I(find_median_inst_mid1_reg[7]), .O(n5368) );
  NR2 U6380 ( .I1(n5368), .I2(find_median_inst_mid2_reg[7]), .O(n5336) );
  INV1S U6381 ( .I(n5336), .O(n5328) );
  ND2S U6382 ( .I1(find_median_inst_mid1_reg[6]), .I2(n5385), .O(n5333) );
  INV1S U6383 ( .I(n5339), .O(n5327) );
  AOI13HS U6384 ( .B1(n5329), .B2(n5328), .B3(n5333), .A1(n5327), .O(n5369) );
  ND2S U6385 ( .I1(find_median_inst_mid3_reg[7]), .I2(n5352), .O(n5330) );
  OR2B1S U6386 ( .I1(n5332), .B1(n5331), .O(n5335) );
  AOI13HS U6387 ( .B1(n5339), .B2(n5338), .B3(n5337), .A1(n5336), .O(n5371) );
  ND2S U6388 ( .I1(find_median_inst_mid3_reg[0]), .I2(n5340), .O(n5342) );
  INV1S U6389 ( .I(find_median_inst_mid3_reg[6]), .O(n5386) );
  ND2S U6390 ( .I1(n5345), .I2(n5344), .O(n5346) );
  MOAI1S U6391 ( .A1(find_median_inst_mid2_reg[6]), .A2(n5386), .B1(n5347), 
        .B2(n5346), .O(n5348) );
  AOI13HS U6392 ( .B1(n5351), .B2(n5350), .B3(n5349), .A1(n5348), .O(n5354) );
  MOAI1S U6393 ( .A1(n5354), .A2(n5353), .B1(find_median_inst_mid3_reg[7]), 
        .B2(n5352), .O(n5355) );
  MOAI1S U6394 ( .A1(n5357), .A2(n5356), .B1(n5371), .B2(n5355), .O(n5389) );
  INV1S U6395 ( .I(find_median_inst_mid3_reg[3]), .O(n5378) );
  FA1S U6396 ( .A(find_median_inst_mid1_reg[1]), .B(
        find_median_inst_mid1_reg[0]), .CI(n5358), .CO(n5359) );
  FA1S U6397 ( .A(n5375), .B(find_median_inst_mid1_reg[2]), .CI(n5359), .CO(
        n5360) );
  ND2S U6398 ( .I1(find_median_inst_mid3_reg[5]), .I2(n5380), .O(n5363) );
  INV1S U6399 ( .I(find_median_inst_mid3_reg[5]), .O(n5381) );
  AOI22S U6400 ( .A1(find_median_inst_mid1_reg[5]), .A2(n5381), .B1(
        find_median_inst_mid1_reg[6]), .B2(n5386), .O(n5365) );
  MOAI1S U6401 ( .A1(find_median_inst_mid1_reg[6]), .A2(n5386), .B1(n5366), 
        .B2(n5365), .O(n5367) );
  INV1S U6402 ( .I(n5370), .O(n5372) );
  AOI22S U6403 ( .A1(n5372), .A2(n5371), .B1(n5370), .B2(n5369), .O(n5382) );
  INV1S U6404 ( .I(n5382), .O(n5388) );
  INV1S U6405 ( .I(n5389), .O(n5384) );
  INV1S U6406 ( .I(n5387), .O(n5390) );
  OAI222S U6407 ( .A1(n5387), .A2(n5375), .B1(n5374), .B2(n5384), .C1(n5373), 
        .C2(n5382), .O(find_median_inst_mid_mid[2]) );
  OAI222S U6408 ( .A1(n5387), .A2(n5378), .B1(n5377), .B2(n5384), .C1(n5376), 
        .C2(n5382), .O(find_median_inst_mid_mid[3]) );
  OAI222S U6409 ( .A1(n5387), .A2(n5381), .B1(n5380), .B2(n5382), .C1(n5379), 
        .C2(n5384), .O(find_median_inst_mid_mid[5]) );
  OAI222S U6410 ( .A1(n5387), .A2(n5386), .B1(n5385), .B2(n5384), .C1(n5383), 
        .C2(n5382), .O(find_median_inst_mid_mid[6]) );
  MOAI1S U6411 ( .A1(n5397), .A2(n5391), .B1(n5397), .B2(
        find_median_inst_min3_reg[1]), .O(find_median_inst_min_max[1]) );
  MOAI1S U6412 ( .A1(n5397), .A2(n5392), .B1(n5397), .B2(
        find_median_inst_min3_reg[2]), .O(find_median_inst_min_max[2]) );
  MOAI1S U6413 ( .A1(n5397), .A2(n5393), .B1(n5397), .B2(
        find_median_inst_min3_reg[3]), .O(find_median_inst_min_max[3]) );
  MOAI1S U6414 ( .A1(n5397), .A2(n5394), .B1(n5397), .B2(
        find_median_inst_min3_reg[4]), .O(find_median_inst_min_max[4]) );
  MOAI1S U6415 ( .A1(n5397), .A2(n5395), .B1(n5397), .B2(
        find_median_inst_min3_reg[5]), .O(find_median_inst_min_max[5]) );
  MOAI1S U6416 ( .A1(n5397), .A2(n5396), .B1(n5397), .B2(
        find_median_inst_min3_reg[6]), .O(find_median_inst_min_max[6]) );
  INV1S U6417 ( .I(find_median_inst_max_min_reg[7]), .O(n5453) );
  NR2 U6418 ( .I1(find_median_inst_mid_mid_reg[7]), .I2(n5453), .O(n5407) );
  INV1S U6419 ( .I(find_median_inst_max_min_reg[6]), .O(n5467) );
  AOI22S U6420 ( .A1(find_median_inst_mid_mid_reg[6]), .A2(n5467), .B1(
        find_median_inst_mid_mid_reg[7]), .B2(n5453), .O(n5406) );
  INV1S U6421 ( .I(find_median_inst_max_min_reg[4]), .O(n5437) );
  INV1S U6422 ( .I(find_median_inst_max_min_reg[5]), .O(n5463) );
  AOI22S U6423 ( .A1(find_median_inst_mid_mid_reg[4]), .A2(n5437), .B1(
        find_median_inst_mid_mid_reg[5]), .B2(n5463), .O(n5404) );
  INV1S U6424 ( .I(find_median_inst_max_min_reg[3]), .O(n5460) );
  INV1S U6425 ( .I(find_median_inst_max_min_reg[2]), .O(n5457) );
  INV1S U6426 ( .I(find_median_inst_max_min_reg[1]), .O(n5430) );
  OAI12HS U6427 ( .B1(find_median_inst_mid_mid_reg[4]), .B2(n5437), .A1(n5400), 
        .O(n5403) );
  INV1S U6428 ( .I(find_median_inst_mid_mid_reg[6]), .O(n5469) );
  INV1S U6429 ( .I(find_median_inst_mid_mid_reg[5]), .O(n5464) );
  AOI22S U6430 ( .A1(find_median_inst_max_min_reg[6]), .A2(n5469), .B1(
        find_median_inst_max_min_reg[5]), .B2(n5464), .O(n5401) );
  OR2B1S U6431 ( .I1(n5407), .B1(n5401), .O(n5402) );
  OAI12HS U6432 ( .B1(n5407), .B2(n5406), .A1(n5405), .O(n5456) );
  INV1S U6433 ( .I(n5456), .O(n5429) );
  INV1S U6434 ( .I(find_median_inst_min_pool_temp[6]), .O(n5470) );
  NR2 U6435 ( .I1(find_median_inst_mid_mid_reg[6]), .I2(n5470), .O(n5422) );
  INV1S U6436 ( .I(find_median_inst_mid_mid_reg[4]), .O(n5410) );
  INV1S U6437 ( .I(find_median_inst_min_pool_temp[5]), .O(n5465) );
  ND2S U6438 ( .I1(n5465), .I2(find_median_inst_mid_mid_reg[5]), .O(n5409) );
  NR2 U6439 ( .I1(n5465), .I2(find_median_inst_mid_mid_reg[5]), .O(n5408) );
  AOI13HS U6440 ( .B1(find_median_inst_min_pool_temp[4]), .B2(n5410), .B3(
        n5409), .A1(n5408), .O(n5421) );
  OA12S U6441 ( .B1(find_median_inst_min_pool_temp[4]), .B2(n5410), .A1(n5409), 
        .O(n5419) );
  INV1S U6442 ( .I(find_median_inst_min_pool_temp[1]), .O(n5431) );
  NR2 U6443 ( .I1(n5431), .I2(find_median_inst_mid_mid_reg[1]), .O(n5413) );
  INV1S U6444 ( .I(find_median_inst_min_pool_temp[2]), .O(n5459) );
  ND2S U6445 ( .I1(find_median_inst_mid_mid_reg[2]), .I2(n5459), .O(n5412) );
  ND2S U6446 ( .I1(find_median_inst_mid_mid_reg[1]), .I2(n5431), .O(n5411) );
  OAI112HS U6447 ( .C1(find_median_inst_min_pool_temp[0]), .C2(n5413), .A1(
        n5412), .B1(n5411), .O(n5416) );
  INV1S U6448 ( .I(find_median_inst_mid_mid_reg[2]), .O(n5458) );
  ND2S U6449 ( .I1(find_median_inst_min_pool_temp[2]), .I2(n5458), .O(n5415)
         );
  INV1S U6450 ( .I(find_median_inst_mid_mid_reg[3]), .O(n5461) );
  ND2S U6451 ( .I1(find_median_inst_min_pool_temp[3]), .I2(n5461), .O(n5414)
         );
  ND3S U6452 ( .I1(n5416), .I2(n5415), .I3(n5414), .O(n5418) );
  INV1S U6453 ( .I(find_median_inst_min_pool_temp[3]), .O(n5462) );
  ND2S U6454 ( .I1(find_median_inst_mid_mid_reg[3]), .I2(n5462), .O(n5417) );
  ND3S U6455 ( .I1(n5419), .I2(n5418), .I3(n5417), .O(n5420) );
  ND2S U6456 ( .I1(find_median_inst_mid_mid_reg[6]), .I2(n5470), .O(n5426) );
  INV1S U6457 ( .I(find_median_inst_min_pool_temp[7]), .O(n5423) );
  ND2S U6458 ( .I1(find_median_inst_mid_mid_reg[7]), .I2(n5423), .O(n5425) );
  NR2 U6459 ( .I1(n5423), .I2(find_median_inst_mid_mid_reg[7]), .O(n5424) );
  AOI13HS U6460 ( .B1(n5427), .B2(n5426), .B3(n5425), .A1(n5424), .O(n5428) );
  MOAI1S U6461 ( .A1(n5429), .A2(n5428), .B1(n5429), .B2(n5428), .O(n5473) );
  AOI22S U6462 ( .A1(find_median_inst_min_pool_temp[6]), .A2(n5467), .B1(
        find_median_inst_min_pool_temp[7]), .B2(n5453), .O(n5451) );
  ND2S U6463 ( .I1(n5465), .I2(find_median_inst_max_min_reg[5]), .O(n5435) );
  NR2 U6464 ( .I1(n5465), .I2(find_median_inst_max_min_reg[5]), .O(n5436) );
  AOI13HS U6465 ( .B1(find_median_inst_min_pool_temp[4]), .B2(n5435), .B3(
        n5437), .A1(n5436), .O(n5446) );
  OA12S U6466 ( .B1(find_median_inst_max_min_reg[3]), .B2(n5462), .A1(n5446), 
        .O(n5450) );
  ND2S U6467 ( .I1(n5457), .I2(find_median_inst_min_pool_temp[2]), .O(n5449)
         );
  INV1S U6468 ( .I(find_median_inst_min_pool_temp[0]), .O(n5432) );
  ND2S U6469 ( .I1(n5430), .I2(find_median_inst_min_pool_temp[1]), .O(n5442)
         );
  MOAI1S U6470 ( .A1(n5457), .A2(find_median_inst_min_pool_temp[2]), .B1(
        find_median_inst_max_min_reg[1]), .B2(n5431), .O(n5441) );
  AO12S U6471 ( .B1(n5432), .B2(n5442), .A1(n5441), .O(n5433) );
  MOAI1S U6472 ( .A1(n5460), .A2(find_median_inst_min_pool_temp[3]), .B1(n5449), .B2(n5433), .O(n5434) );
  ND2S U6473 ( .I1(n5450), .I2(n5434), .O(n5439) );
  OA13S U6474 ( .B1(n5437), .B2(n5436), .B3(find_median_inst_min_pool_temp[4]), 
        .A1(n5435), .O(n5444) );
  ND2S U6475 ( .I1(find_median_inst_max_min_reg[6]), .I2(n5470), .O(n5438) );
  MOAI1S U6476 ( .A1(find_median_inst_min_pool_temp[7]), .A2(n5453), .B1(n5451), .B2(n5440), .O(n5455) );
  AO12S U6477 ( .B1(find_median_inst_max_min_reg[0]), .B2(n5442), .A1(n5441), 
        .O(n5448) );
  ND2S U6478 ( .I1(find_median_inst_max_min_reg[3]), .I2(n5462), .O(n5443) );
  ND2S U6479 ( .I1(n5444), .I2(n5443), .O(n5445) );
  MOAI1S U6480 ( .A1(find_median_inst_min_pool_temp[6]), .A2(n5467), .B1(n5446), .B2(n5445), .O(n5447) );
  AO13S U6481 ( .B1(n5450), .B2(n5449), .B3(n5448), .A1(n5447), .O(n5452) );
  MOAI1S U6482 ( .A1(n5453), .A2(find_median_inst_min_pool_temp[7]), .B1(n5452), .B2(n5451), .O(n5454) );
  MOAI1S U6483 ( .A1(n5456), .A2(n5455), .B1(n5456), .B2(n5454), .O(n5472) );
  INV1S U6484 ( .I(n5472), .O(n5466) );
  INV1S U6485 ( .I(n5473), .O(n5468) );
  INV1S U6486 ( .I(n5471), .O(n5474) );
  OAI222S U6487 ( .A1(n5471), .A2(n5459), .B1(n5458), .B2(n5468), .C1(n5457), 
        .C2(n5466), .O(find_median_inst_final_mid[2]) );
  OAI222S U6488 ( .A1(n5471), .A2(n5462), .B1(n5461), .B2(n5468), .C1(n5460), 
        .C2(n5466), .O(find_median_inst_final_mid[3]) );
  OAI222S U6489 ( .A1(n5471), .A2(n5465), .B1(n5464), .B2(n5468), .C1(n5463), 
        .C2(n5466), .O(find_median_inst_final_mid[5]) );
  OAI222S U6490 ( .A1(n5471), .A2(n5470), .B1(n5469), .B2(n5468), .C1(n5467), 
        .C2(n5466), .O(find_median_inst_final_mid[6]) );
  ND2S U6491 ( .I1(median_in[53]), .I2(n5913), .O(n5476) );
  MOAI1S U6492 ( .A1(n5913), .A2(median_in[53]), .B1(n5926), .B2(median_in[70]), .O(n5475) );
  AOI13HS U6493 ( .B1(median_in[68]), .B2(n5904), .B3(n5476), .A1(n5475), .O(
        n5484) );
  AOI22S U6494 ( .A1(median_in[53]), .A2(n5913), .B1(median_in[52]), .B2(n5532), .O(n5479) );
  ND2S U6495 ( .I1(n5480), .I2(n5479), .O(n5483) );
  ND2S U6496 ( .I1(median_in[54]), .I2(n5927), .O(n5481) );
  NR2 U6497 ( .I1(median_in[65]), .I2(n5525), .O(n5486) );
  OAI12HS U6498 ( .B1(n5486), .B2(median_in[56]), .A1(n5485), .O(n5488) );
  ND2S U6499 ( .I1(n5488), .I2(n5487), .O(n5489) );
  ND3S U6500 ( .I1(n5491), .I2(n5490), .I3(n5489), .O(n5493) );
  AOI13HS U6501 ( .B1(n5495), .B2(n5494), .B3(n5493), .A1(n5492), .O(n5497) );
  OAI22S U6502 ( .A1(n5497), .A2(n5496), .B1(n5945), .B2(median_in[63]), .O(
        n5503) );
  INV1S U6503 ( .I(n5502), .O(n5498) );
  NR2 U6504 ( .I1(n5499), .I2(n5498), .O(n5500) );
  NR2 U6505 ( .I1(n5503), .I2(n5500), .O(n5501) );
  AOI13HS U6506 ( .B1(n5520), .B2(n5542), .B3(n5502), .A1(n5501), .O(n5529) );
  INV1S U6507 ( .I(n5503), .O(n5523) );
  INV1S U6508 ( .I(n5504), .O(n5505) );
  OAI12HS U6509 ( .B1(median_in[54]), .B2(n5928), .A1(n5505), .O(n5518) );
  AOI22S U6510 ( .A1(median_in[51]), .A2(n5895), .B1(median_in[50]), .B2(n5527), .O(n5510) );
  NR2 U6511 ( .I1(median_in[57]), .I2(n5526), .O(n5508) );
  ND2S U6512 ( .I1(median_in[58]), .I2(n5528), .O(n5507) );
  MOAI1S U6513 ( .A1(median_in[49]), .A2(n5525), .B1(n5528), .B2(median_in[58]), .O(n5506) );
  MAOI1S U6514 ( .A1(n5508), .A2(n5507), .B1(n6320), .B2(n5506), .O(n5509) );
  AOI22S U6515 ( .A1(median_in[59]), .A2(n5893), .B1(n5510), .B2(n5509), .O(
        n5517) );
  NR2 U6516 ( .I1(median_in[62]), .I2(n5926), .O(n5515) );
  OR2S U6517 ( .I1(median_in[60]), .I2(n5904), .O(n5511) );
  ND2S U6518 ( .I1(median_in[53]), .I2(n5914), .O(n5513) );
  OR3B2S U6519 ( .I1(n5515), .B1(n5511), .B2(n5513), .O(n5516) );
  NR2 U6520 ( .I1(median_in[53]), .I2(n5914), .O(n5512) );
  AOI13HS U6521 ( .B1(median_in[60]), .B2(n5904), .B3(n5513), .A1(n5512), .O(
        n5514) );
  OAI22S U6522 ( .A1(n5517), .A2(n5516), .B1(n5515), .B2(n5514), .O(n5519) );
  OAI12HS U6523 ( .B1(n5518), .B2(n5519), .A1(n5540), .O(n5522) );
  AOI22S U6524 ( .A1(n5523), .A2(n5522), .B1(n5521), .B2(n5520), .O(n5530) );
  OAI222S U6525 ( .A1(n5531), .A2(n6320), .B1(n5545), .B2(n5529), .C1(n5524), 
        .C2(n5530), .O(find_median_inst_mid1[0]) );
  OAI222S U6526 ( .A1(n5531), .A2(n5526), .B1(n5525), .B2(n5530), .C1(n5534), 
        .C2(n5529), .O(find_median_inst_mid1[1]) );
  OAI222S U6527 ( .A1(n5531), .A2(n5528), .B1(n5527), .B2(n5530), .C1(n5533), 
        .C2(n5529), .O(find_median_inst_mid1[2]) );
  OAI222S U6528 ( .A1(n5531), .A2(n5893), .B1(n5895), .B2(n5530), .C1(n5894), 
        .C2(n5529), .O(find_median_inst_mid1[3]) );
  OAI222S U6529 ( .A1(n5531), .A2(n5904), .B1(n5902), .B2(n5530), .C1(n5532), 
        .C2(n5529), .O(find_median_inst_mid1[4]) );
  OAI222S U6530 ( .A1(n5531), .A2(n6321), .B1(n5914), .B2(n5530), .C1(n5913), 
        .C2(n5529), .O(find_median_inst_mid1[5]) );
  OAI222S U6531 ( .A1(n5531), .A2(n5926), .B1(n5927), .B2(n5529), .C1(n5928), 
        .C2(n5530), .O(find_median_inst_mid1[6]) );
  OAI222S U6532 ( .A1(n5531), .A2(n5940), .B1(n5944), .B2(n5530), .C1(n5945), 
        .C2(n5529), .O(find_median_inst_mid1[7]) );
  MOAI1S U6533 ( .A1(n5546), .A2(median_in[62]), .B1(n5546), .B2(n5927), .O(
        n5553) );
  MOAI1S U6534 ( .A1(n5546), .A2(median_in[61]), .B1(n5546), .B2(n5913), .O(
        n5552) );
  MOAI1S U6535 ( .A1(n5546), .A2(median_in[60]), .B1(n5546), .B2(n5532), .O(
        n5551) );
  MOAI1S U6536 ( .A1(n5546), .A2(median_in[59]), .B1(n5546), .B2(n5894), .O(
        n5550) );
  MOAI1S U6537 ( .A1(n5546), .A2(median_in[58]), .B1(n5546), .B2(n5533), .O(
        n5549) );
  FA1S U6538 ( .A(median_in[49]), .B(median_in[48]), .CI(n5548), .CO(n5535) );
  FA1S U6539 ( .A(n5549), .B(median_in[50]), .CI(n5535), .CO(n5536) );
  FA1S U6540 ( .A(n5550), .B(median_in[51]), .CI(n5536), .CO(n5537) );
  FA1S U6541 ( .A(median_in[52]), .B(n5551), .CI(n5537), .CO(n5538) );
  MOAI1S U6542 ( .A1(n5546), .A2(median_in[56]), .B1(n5546), .B2(n5545), .O(
        n5547) );
  MOAI1S U6543 ( .A1(n5554), .A2(n5547), .B1(n5554), .B2(median_in[48]), .O(
        find_median_inst_min1[0]) );
  MOAI1S U6544 ( .A1(n5554), .A2(n5548), .B1(n5554), .B2(median_in[49]), .O(
        find_median_inst_min1[1]) );
  MOAI1S U6545 ( .A1(n5554), .A2(n5549), .B1(n5554), .B2(median_in[50]), .O(
        find_median_inst_min1[2]) );
  MOAI1S U6546 ( .A1(n5554), .A2(n5550), .B1(n5554), .B2(median_in[51]), .O(
        find_median_inst_min1[3]) );
  MOAI1S U6547 ( .A1(n5554), .A2(n5551), .B1(n5554), .B2(median_in[52]), .O(
        find_median_inst_min1[4]) );
  MOAI1S U6548 ( .A1(n5554), .A2(n5552), .B1(n5554), .B2(median_in[53]), .O(
        find_median_inst_min1[5]) );
  MOAI1S U6549 ( .A1(n5554), .A2(n5553), .B1(n5554), .B2(median_in[54]), .O(
        find_median_inst_min1[6]) );
  NR3 U6550 ( .I1(n5945), .I2(n5940), .I3(n5944), .O(find_median_inst_min1[7])
         );
  MOAI1S U6551 ( .A1(n5556), .A2(n5555), .B1(n5556), .B2(median_in[54]), .O(
        find_median_inst_max1[6]) );
  INV1S U6552 ( .I(SRAM_64X32_WE), .O(n3416) );
  INV1S U6553 ( .I(SRAM_192X32_WE), .O(n3415) );
  OAI12HS U6554 ( .B1(n5558), .B2(n3517), .A1(n5557), .O(n3401) );
  MOAI1S U6555 ( .A1(set_count[0]), .A2(n5591), .B1(set_count[0]), .B2(n5559), 
        .O(n3400) );
  INV1S U6556 ( .I(set_count[2]), .O(n5563) );
  NR2 U6557 ( .I1(set_count[0]), .I2(n5591), .O(n5560) );
  NR2 U6558 ( .I1(n5560), .I2(n5559), .O(n5719) );
  OA12S U6559 ( .B1(set_count[1]), .B2(n5591), .A1(n5719), .O(n5562) );
  MOAI1S U6560 ( .A1(n5563), .A2(n5562), .B1(n5563), .B2(n5561), .O(n3399) );
  NR2 U6561 ( .I1(action_idx[0]), .I2(in_valid2), .O(n5564) );
  NR2 U6562 ( .I1(n5565), .I2(n5564), .O(n3398) );
  AOI22S U6563 ( .A1(action_idx[1]), .A2(n5565), .B1(n5566), .B2(n5576), .O(
        n3397) );
  NR2 U6564 ( .I1(n5576), .I2(n5566), .O(n5579) );
  NR2 U6565 ( .I1(action_idx[3]), .I2(n5568), .O(n5570) );
  INV1S U6566 ( .I(n5570), .O(n5571) );
  INV1S U6567 ( .I(action[0]), .O(n5586) );
  MOAI1S U6568 ( .A1(n5571), .A2(n5586), .B1(n5571), .B2(action_reg_7__0_), 
        .O(n3394) );
  INV1S U6569 ( .I(action[2]), .O(n5587) );
  MOAI1S U6570 ( .A1(n5571), .A2(n5587), .B1(n5571), .B2(action_reg_7__2_), 
        .O(n3393) );
  INV1S U6571 ( .I(action[1]), .O(n5588) );
  MOAI1S U6572 ( .A1(n5571), .A2(n5588), .B1(n5571), .B2(action_reg_7__1_), 
        .O(n3392) );
  OR2B1S U6573 ( .I1(action_idx[3]), .B1(action_idx[2]), .O(n5574) );
  NR3 U6574 ( .I1(action_idx[0]), .I2(n5572), .I3(n5574), .O(n5577) );
  MOAI1S U6575 ( .A1(n5573), .A2(n5586), .B1(n5573), .B2(action_reg_6__0_), 
        .O(n3391) );
  MOAI1S U6576 ( .A1(n5573), .A2(n5587), .B1(n5573), .B2(action_reg_6__2_), 
        .O(n3390) );
  MOAI1S U6577 ( .A1(n5573), .A2(n5588), .B1(n5573), .B2(action_reg_6__1_), 
        .O(n3389) );
  ND3S U6578 ( .I1(action_idx[0]), .I2(in_valid2), .I3(n5576), .O(n5584) );
  MOAI1S U6579 ( .A1(n5575), .A2(n5586), .B1(n5575), .B2(action_reg_5__0_), 
        .O(n3388) );
  MOAI1S U6580 ( .A1(n5575), .A2(n5587), .B1(n5575), .B2(action_reg_5__2_), 
        .O(n3387) );
  MOAI1S U6581 ( .A1(n5575), .A2(n5588), .B1(n5575), .B2(action_reg_5__1_), 
        .O(n3386) );
  MOAI1S U6582 ( .A1(n5578), .A2(n5586), .B1(n5578), .B2(action_reg_4__0_), 
        .O(n3385) );
  MOAI1S U6583 ( .A1(n5578), .A2(n5587), .B1(n5578), .B2(action_reg_4__2_), 
        .O(n3384) );
  MOAI1S U6584 ( .A1(n5578), .A2(n5588), .B1(n5578), .B2(action_reg_4__1_), 
        .O(n3383) );
  MOAI1S U6585 ( .A1(n5581), .A2(n5586), .B1(n5581), .B2(action_reg_3__0_), 
        .O(n3382) );
  MOAI1S U6586 ( .A1(n5581), .A2(n5587), .B1(n5581), .B2(action_reg_3__2_), 
        .O(n3381) );
  MOAI1S U6587 ( .A1(n5581), .A2(n5588), .B1(n5581), .B2(action_reg_3__1_), 
        .O(n3380) );
  MOAI1S U6588 ( .A1(n5583), .A2(n5586), .B1(n5583), .B2(action_reg_2__0_), 
        .O(n3379) );
  MOAI1S U6589 ( .A1(n5583), .A2(n5587), .B1(n5583), .B2(action_reg_2__2_), 
        .O(n3378) );
  MOAI1S U6590 ( .A1(n5583), .A2(n5588), .B1(n5583), .B2(action_reg_2__1_), 
        .O(n3377) );
  MOAI1S U6591 ( .A1(n5589), .A2(n5586), .B1(n5589), .B2(action_reg_1__0_), 
        .O(n3376) );
  MOAI1S U6592 ( .A1(n5589), .A2(n5587), .B1(n5589), .B2(action_reg_1__2_), 
        .O(n3375) );
  MOAI1S U6593 ( .A1(n5589), .A2(n5588), .B1(n5589), .B2(action_reg_1__1_), 
        .O(n3374) );
  AN2S U6594 ( .I1(n5590), .I2(n5591), .O(n3371) );
  ND2S U6595 ( .I1(conv_dly3[0]), .I2(conv_dly3[1]), .O(n5592) );
  OAI22S U6596 ( .A1(n5600), .A2(n5594), .B1(n3517), .B2(n5593), .O(n3370) );
  INV1S U6597 ( .I(conv_dly3[0]), .O(n5597) );
  OAI12HS U6598 ( .B1(conv_dly3[1]), .B2(n5594), .A1(n5597), .O(n5595) );
  AOI22S U6599 ( .A1(n3517), .A2(n5597), .B1(n5596), .B2(n5595), .O(n3369) );
  NR2 U6600 ( .I1(n3517), .I2(n5597), .O(n5598) );
  NR2 U6601 ( .I1(conv_dly3[1]), .I2(n5598), .O(n5599) );
  NR2 U6602 ( .I1(n5600), .I2(n5599), .O(n3368) );
  MOAI1S U6603 ( .A1(n5601), .A2(n5608), .B1(n5607), .B2(max_temp[0]), .O(
        n3361) );
  MOAI1S U6604 ( .A1(n5602), .A2(n5608), .B1(max_temp[1]), .B2(n5607), .O(
        n3360) );
  MOAI1S U6605 ( .A1(n5603), .A2(n5608), .B1(max_temp[2]), .B2(n5607), .O(
        n3359) );
  MOAI1S U6606 ( .A1(n5604), .A2(n5608), .B1(max_temp[3]), .B2(n5607), .O(
        n3358) );
  MOAI1S U6607 ( .A1(n5605), .A2(n5608), .B1(max_temp[4]), .B2(n5607), .O(
        n3357) );
  MOAI1S U6608 ( .A1(n5606), .A2(n5608), .B1(max_temp[5]), .B2(n5607), .O(
        n3356) );
  MOAI1S U6609 ( .A1(n5609), .A2(n5608), .B1(max_temp[7]), .B2(n5607), .O(
        n3355) );
  NR2 U6610 ( .I1(n5610), .I2(n5626), .O(n5621) );
  FA1S U6611 ( .A(image[3]), .B(wgt_temp[2]), .CI(n5614), .CO(n5616), .S(n5615) );
  FA1S U6612 ( .A(image[5]), .B(wgt_temp[4]), .CI(n5618), .CO(n5620), .S(n5619) );
  FA1S U6613 ( .A(image[7]), .B(wgt_temp[6]), .CI(n5623), .CO(n3674), .S(n5625) );
  ND2S U6614 ( .I1(n3493), .I2(template_count[3]), .O(n5628) );
  MOAI1S U6615 ( .A1(n5631), .A2(n5628), .B1(n5631), .B2(n5627), .O(n3346) );
  NR2 U6616 ( .I1(template_count[2]), .I2(n5629), .O(n5630) );
  NR3 U6617 ( .I1(n5631), .I2(n3492), .I3(n5630), .O(n3345) );
  AOI22S U6618 ( .A1(n5636), .A2(n5633), .B1(template_count[1]), .B2(n5632), 
        .O(n5634) );
  NR2 U6619 ( .I1(n5634), .I2(n3492), .O(n3344) );
  MOAI1S U6620 ( .A1(template_count[0]), .A2(n3492), .B1(n5636), .B2(n5635), 
        .O(n3343) );
  INV1S U6621 ( .I(template[7]), .O(n5645) );
  MOAI1S U6622 ( .A1(n5637), .A2(n5645), .B1(n5637), .B2(template_reg[7]), .O(
        n3341) );
  INV1S U6623 ( .I(template[6]), .O(n5646) );
  MOAI1S U6624 ( .A1(n5637), .A2(n5646), .B1(n5637), .B2(template_reg[6]), .O(
        n3340) );
  INV1S U6625 ( .I(template[5]), .O(n5647) );
  MOAI1S U6626 ( .A1(n5637), .A2(n5647), .B1(n5637), .B2(template_reg[5]), .O(
        n3339) );
  MOAI1S U6627 ( .A1(n5638), .A2(n5645), .B1(n5638), .B2(template_reg[15]), 
        .O(n3333) );
  MOAI1S U6628 ( .A1(n5638), .A2(n5646), .B1(n5638), .B2(template_reg[14]), 
        .O(n3332) );
  MOAI1S U6629 ( .A1(n5638), .A2(n5647), .B1(n5638), .B2(template_reg[13]), 
        .O(n3331) );
  MOAI1S U6630 ( .A1(n5639), .A2(n5645), .B1(n5639), .B2(template_reg[23]), 
        .O(n3325) );
  MOAI1S U6631 ( .A1(n5639), .A2(n5646), .B1(n5639), .B2(template_reg[22]), 
        .O(n3324) );
  MOAI1S U6632 ( .A1(n5639), .A2(n5647), .B1(n5639), .B2(template_reg[21]), 
        .O(n3323) );
  MOAI1S U6633 ( .A1(n5640), .A2(n5645), .B1(n5640), .B2(template_reg[31]), 
        .O(n3317) );
  MOAI1S U6634 ( .A1(n5640), .A2(n5646), .B1(n5640), .B2(template_reg[30]), 
        .O(n3316) );
  MOAI1S U6635 ( .A1(n5640), .A2(n5647), .B1(n5640), .B2(template_reg[29]), 
        .O(n3315) );
  MOAI1S U6636 ( .A1(n5641), .A2(n5645), .B1(n5641), .B2(template_reg[39]), 
        .O(n3309) );
  MOAI1S U6637 ( .A1(n5641), .A2(n5646), .B1(n5641), .B2(template_reg[38]), 
        .O(n3308) );
  MOAI1S U6638 ( .A1(n5641), .A2(n5647), .B1(n5641), .B2(template_reg[37]), 
        .O(n3307) );
  MOAI1S U6639 ( .A1(n5642), .A2(n5645), .B1(n5642), .B2(template_reg[47]), 
        .O(n3301) );
  MOAI1S U6640 ( .A1(n5642), .A2(n5646), .B1(n5642), .B2(template_reg[46]), 
        .O(n3300) );
  MOAI1S U6641 ( .A1(n5642), .A2(n5647), .B1(n5642), .B2(template_reg[45]), 
        .O(n3299) );
  MOAI1S U6642 ( .A1(n5643), .A2(n5645), .B1(n5643), .B2(template_reg[55]), 
        .O(n3293) );
  MOAI1S U6643 ( .A1(n5643), .A2(n5646), .B1(n5643), .B2(template_reg[54]), 
        .O(n3292) );
  MOAI1S U6644 ( .A1(n5643), .A2(n5647), .B1(n5643), .B2(template_reg[53]), 
        .O(n3291) );
  MOAI1S U6645 ( .A1(n5644), .A2(n5645), .B1(n5644), .B2(template_reg[63]), 
        .O(n3285) );
  MOAI1S U6646 ( .A1(n5644), .A2(n5646), .B1(n5644), .B2(template_reg[62]), 
        .O(n3284) );
  MOAI1S U6647 ( .A1(n5644), .A2(n5647), .B1(n5644), .B2(template_reg[61]), 
        .O(n3283) );
  MOAI1S U6648 ( .A1(n61240), .A2(n5645), .B1(n61240), .B2(template_reg[71]), 
        .O(n3277) );
  MOAI1S U6649 ( .A1(n61240), .A2(n5646), .B1(n61240), .B2(template_reg[70]), 
        .O(n3276) );
  MOAI1S U6650 ( .A1(n61240), .A2(n5647), .B1(n61240), .B2(template_reg[69]), 
        .O(n3275) );
  INV1S U6651 ( .I(SRAM_192_32_in_count[0]), .O(n5651) );
  NR2 U6652 ( .I1(n5651), .I2(n5650), .O(n5653) );
  OAI22S U6653 ( .A1(SRAM_192_32_in_count[1]), .A2(n5653), .B1(n5648), .B2(
        n5650), .O(n5649) );
  NR2 U6654 ( .I1(n5654), .I2(n5649), .O(n3270) );
  AN2S U6655 ( .I1(n5651), .I2(n5650), .O(n5652) );
  NR3 U6656 ( .I1(n5654), .I2(n5653), .I3(n5652), .O(n3269) );
  ND2S U6657 ( .I1(n5656), .I2(n5655), .O(n5658) );
  OAI22S U6658 ( .A1(n5709), .A2(n5658), .B1(n5657), .B2(n5656), .O(n3235) );
  MOAI1S U6659 ( .A1(n5659), .A2(n3488), .B1(n5659), .B2(n3488), .O(n5660) );
  MOAI1S U6660 ( .A1(n3488), .A2(n6301), .B1(n5715), .B2(n5660), .O(n3233) );
  MOAI1S U6661 ( .A1(current_action_idx[0]), .A2(n5665), .B1(
        current_action_idx[0]), .B2(n5661), .O(n3232) );
  ND2S U6662 ( .I1(n5662), .I2(current_action_idx[0]), .O(n5664) );
  OAI22S U6663 ( .A1(n5665), .A2(n5664), .B1(n5663), .B2(n5662), .O(n3231) );
  NR2 U6664 ( .I1(n5725), .I2(n5678), .O(n5671) );
  INV1S U6665 ( .I(n5671), .O(n5666) );
  OAI112HS U6666 ( .C1(n61230), .C2(n5668), .A1(n5667), .B1(n5666), .O(n3229)
         );
  ND2S U6667 ( .I1(n5670), .I2(n5669), .O(n5674) );
  NR2 U6668 ( .I1(n5672), .I2(n5671), .O(n5673) );
  ND3S U6669 ( .I1(n5674), .I2(n5673), .I3(n5675), .O(n5676) );
  OAI22S U6670 ( .A1(n61230), .A2(n5676), .B1(n5675), .B2(n5674), .O(n3228) );
  INV1S U6671 ( .I(n5677), .O(n5684) );
  ND2S U6672 ( .I1(n5678), .I2(n5684), .O(n5681) );
  OAI222S U6673 ( .A1(n5680), .A2(n5679), .B1(n5681), .B2(n6309), .C1(n61250), 
        .C2(n5684), .O(n3227) );
  INV1S U6674 ( .I(image_size_reg[1]), .O(n61260) );
  ND2S U6675 ( .I1(n5682), .I2(n5681), .O(n5683) );
  MOAI1S U6676 ( .A1(n5684), .A2(n61260), .B1(image_size_temp[1]), .B2(n5683), 
        .O(n3226) );
  MOAI1S U6677 ( .A1(cal_count[5]), .A2(n5687), .B1(cal_count[5]), .B2(n5687), 
        .O(n5685) );
  MOAI1S U6678 ( .A1(n5686), .A2(n6301), .B1(n5715), .B2(n5685), .O(n3225) );
  ND2S U6679 ( .I1(n5688), .I2(n5687), .O(n5689) );
  MOAI1S U6680 ( .A1(n5709), .A2(n5689), .B1(cal_count[4]), .B2(n5695), .O(
        n3224) );
  NR2 U6681 ( .I1(n5727), .I2(n5728), .O(n5691) );
  OAI22S U6682 ( .A1(n5691), .A2(n5709), .B1(n5690), .B2(n6301), .O(n3221) );
  MOAI1S U6683 ( .A1(n5692), .A2(n6301), .B1(n5692), .B2(n5715), .O(n3220) );
  ND3S U6684 ( .I1(cal_count_10[2]), .I2(n5693), .I3(n6301), .O(n5700) );
  INV1S U6685 ( .I(cal_count_10[3]), .O(n5699) );
  ND2S U6686 ( .I1(n5699), .I2(n5712), .O(n5698) );
  NR2 U6687 ( .I1(cal_count_10[0]), .I2(n5709), .O(n5694) );
  NR2 U6688 ( .I1(n5695), .I2(n5694), .O(n5707) );
  AOI22S U6689 ( .A1(n5700), .A2(n5699), .B1(n5698), .B2(n5702), .O(n3219) );
  OAI22S U6690 ( .A1(n5703), .A2(n5702), .B1(n5709), .B2(n5701), .O(n3218) );
  NR2 U6691 ( .I1(n5705), .I2(n5704), .O(n5706) );
  MOAI1S U6692 ( .A1(n5708), .A2(n5707), .B1(n5708), .B2(n5706), .O(n3216) );
  MOAI1S U6693 ( .A1(n5710), .A2(n5709), .B1(cal_count_5[1]), .B2(n5711), .O(
        n3214) );
  AOI13HS U6694 ( .B1(n5714), .B2(n5713), .B3(n5712), .A1(n5711), .O(n5716) );
  MOAI1S U6695 ( .A1(n5716), .A2(n6024), .B1(n5984), .B2(n5715), .O(n3213) );
  AOI22S U6696 ( .A1(set_count[1]), .A2(n5719), .B1(n5718), .B2(n5717), .O(
        n3197) );
  AOI22S U6697 ( .A1(n5725), .A2(n6244), .B1(n5766), .B2(n5724), .O(n5726) );
  NR2 U6698 ( .I1(n5726), .I2(n6245), .O(n5730) );
  INV1S U6699 ( .I(median_result[0]), .O(n5731) );
  MOAI1S U6700 ( .A1(n5738), .A2(n5731), .B1(n5738), .B2(filter_result_reg[64]), .O(n3195) );
  MOAI1S U6701 ( .A1(n5739), .A2(n5731), .B1(n5739), .B2(filter_result_reg[72]), .O(n3194) );
  MOAI1S U6702 ( .A1(n5740), .A2(n5731), .B1(n5740), .B2(filter_result_reg[80]), .O(n3193) );
  MOAI1S U6703 ( .A1(n5742), .A2(n5731), .B1(n5742), .B2(filter_result_reg[88]), .O(n3192) );
  INV1S U6704 ( .I(median_result[1]), .O(n5732) );
  MOAI1S U6705 ( .A1(n5738), .A2(n5732), .B1(n5738), .B2(filter_result_reg[65]), .O(n3191) );
  MOAI1S U6706 ( .A1(n5739), .A2(n5732), .B1(n5739), .B2(filter_result_reg[73]), .O(n3190) );
  MOAI1S U6707 ( .A1(n5740), .A2(n5732), .B1(n5740), .B2(filter_result_reg[81]), .O(n3189) );
  MOAI1S U6708 ( .A1(n5742), .A2(n5732), .B1(n5742), .B2(filter_result_reg[89]), .O(n3188) );
  INV1S U6709 ( .I(median_result[2]), .O(n5733) );
  MOAI1S U6710 ( .A1(n5738), .A2(n5733), .B1(n5738), .B2(filter_result_reg[66]), .O(n3187) );
  MOAI1S U6711 ( .A1(n5739), .A2(n5733), .B1(n5739), .B2(filter_result_reg[74]), .O(n3186) );
  MOAI1S U6712 ( .A1(n5740), .A2(n5733), .B1(n5740), .B2(filter_result_reg[82]), .O(n3185) );
  MOAI1S U6713 ( .A1(n5742), .A2(n5733), .B1(n5742), .B2(filter_result_reg[90]), .O(n3184) );
  INV1S U6714 ( .I(median_result[3]), .O(n5734) );
  MOAI1S U6715 ( .A1(n5738), .A2(n5734), .B1(n5738), .B2(filter_result_reg[67]), .O(n3183) );
  MOAI1S U6716 ( .A1(n5739), .A2(n5734), .B1(n5739), .B2(filter_result_reg[75]), .O(n3182) );
  MOAI1S U6717 ( .A1(n5740), .A2(n5734), .B1(n5740), .B2(filter_result_reg[83]), .O(n3181) );
  MOAI1S U6718 ( .A1(n5742), .A2(n5734), .B1(n5742), .B2(filter_result_reg[91]), .O(n3180) );
  INV1S U6719 ( .I(median_result[4]), .O(n5735) );
  MOAI1S U6720 ( .A1(n5738), .A2(n5735), .B1(n5738), .B2(filter_result_reg[68]), .O(n3179) );
  MOAI1S U6721 ( .A1(n5739), .A2(n5735), .B1(n5739), .B2(filter_result_reg[76]), .O(n3178) );
  MOAI1S U6722 ( .A1(n5740), .A2(n5735), .B1(n5740), .B2(filter_result_reg[84]), .O(n3177) );
  MOAI1S U6723 ( .A1(n5742), .A2(n5735), .B1(n5742), .B2(filter_result_reg[92]), .O(n3176) );
  INV1S U6724 ( .I(median_result[5]), .O(n5736) );
  MOAI1S U6725 ( .A1(n5738), .A2(n5736), .B1(n5738), .B2(filter_result_reg[69]), .O(n3175) );
  MOAI1S U6726 ( .A1(n5739), .A2(n5736), .B1(n5739), .B2(filter_result_reg[77]), .O(n3174) );
  MOAI1S U6727 ( .A1(n5740), .A2(n5736), .B1(n5740), .B2(filter_result_reg[85]), .O(n3173) );
  MOAI1S U6728 ( .A1(n5742), .A2(n5736), .B1(n5742), .B2(filter_result_reg[93]), .O(n3172) );
  INV1S U6729 ( .I(median_result[6]), .O(n5737) );
  MOAI1S U6730 ( .A1(n5738), .A2(n5737), .B1(n5738), .B2(filter_result_reg[70]), .O(n3171) );
  MOAI1S U6731 ( .A1(n5739), .A2(n5737), .B1(n5739), .B2(filter_result_reg[78]), .O(n3170) );
  MOAI1S U6732 ( .A1(n5740), .A2(n5737), .B1(n5740), .B2(filter_result_reg[86]), .O(n3169) );
  MOAI1S U6733 ( .A1(n5742), .A2(n5737), .B1(n5742), .B2(filter_result_reg[94]), .O(n3168) );
  INV1S U6734 ( .I(median_result[7]), .O(n5741) );
  MOAI1S U6735 ( .A1(n5738), .A2(n5741), .B1(n5738), .B2(filter_result_reg[71]), .O(n3167) );
  MOAI1S U6736 ( .A1(n5739), .A2(n5741), .B1(n5739), .B2(filter_result_reg[79]), .O(n3166) );
  MOAI1S U6737 ( .A1(n5740), .A2(n5741), .B1(n5740), .B2(filter_result_reg[87]), .O(n3165) );
  MOAI1S U6738 ( .A1(n5742), .A2(n5741), .B1(n5742), .B2(filter_result_reg[95]), .O(n3164) );
  AN2 U6739 ( .I1(n5744), .I2(n5743), .O(n6056) );
  MOAI1S U6740 ( .A1(n5933), .A2(n5861), .B1(n5933), .B2(SRAM_out_buffer[32]), 
        .O(n3162) );
  MOAI1S U6741 ( .A1(n5934), .A2(n5861), .B1(n5934), .B2(SRAM_out_buffer[64]), 
        .O(n3161) );
  NR2 U6742 ( .I1(n5746), .I2(n5745), .O(n5747) );
  MOAI1S U6743 ( .A1(n5750), .A2(n5749), .B1(n5748), .B2(n5747), .O(n5754) );
  OAI22S U6744 ( .A1(n5752), .A2(n3486), .B1(n5751), .B2(n5754), .O(n5762) );
  AOI22S U6745 ( .A1(n5755), .A2(n5754), .B1(n5753), .B2(n5752), .O(n5757) );
  AOI13HS U6746 ( .B1(n5764), .B2(n5761), .B3(n5760), .A1(n5759), .O(n6057) );
  OAI12HS U6747 ( .B1(n5763), .B2(n5762), .A1(n6057), .O(n6060) );
  INV1S U6748 ( .I(n6057), .O(n5932) );
  NR2 U6749 ( .I1(n5764), .I2(n6245), .O(n5930) );
  MOAI1S U6750 ( .A1(n5933), .A2(n5867), .B1(n5933), .B2(SRAM_out_buffer[34]), 
        .O(n3156) );
  MOAI1S U6751 ( .A1(n5933), .A2(n5870), .B1(n5933), .B2(SRAM_out_buffer[35]), 
        .O(n3153) );
  INV1S U6752 ( .I(n5793), .O(n5873) );
  MOAI1S U6753 ( .A1(n5933), .A2(n5873), .B1(n5933), .B2(SRAM_out_buffer[36]), 
        .O(n3150) );
  MOAI1S U6754 ( .A1(n5934), .A2(n5873), .B1(n5934), .B2(SRAM_out_buffer[68]), 
        .O(n3149) );
  MOAI1S U6755 ( .A1(n5934), .A2(n5876), .B1(n5934), .B2(SRAM_out_buffer[69]), 
        .O(n3146) );
  MOAI1S U6756 ( .A1(n5934), .A2(n5881), .B1(n5934), .B2(SRAM_out_buffer[70]), 
        .O(n3143) );
  INV1S U6757 ( .I(n5850), .O(n5858) );
  MOAI1S U6758 ( .A1(n5933), .A2(n5858), .B1(n5933), .B2(SRAM_out_buffer[39]), 
        .O(n3141) );
  MOAI1S U6759 ( .A1(n5934), .A2(n5858), .B1(n5934), .B2(SRAM_out_buffer[71]), 
        .O(n3140) );
  MOAI1S U6760 ( .A1(n5934), .A2(n5860), .B1(n5934), .B2(SRAM_out_buffer[72]), 
        .O(n3137) );
  ND3S U6761 ( .I1(n6243), .I2(n5767), .I3(n5766), .O(n5768) );
  INV1S U6762 ( .I(n5930), .O(n6062) );
  INV1S U6763 ( .I(n6062), .O(n5916) );
  MOAI1S U6764 ( .A1(n5934), .A2(n5863), .B1(n5934), .B2(SRAM_out_buffer[73]), 
        .O(n3131) );
  MOAI1S U6765 ( .A1(n5934), .A2(n5866), .B1(n5934), .B2(SRAM_out_buffer[74]), 
        .O(n3125) );
  MOAI1S U6766 ( .A1(n5934), .A2(n5869), .B1(n5934), .B2(SRAM_out_buffer[75]), 
        .O(n3119) );
  MOAI1S U6767 ( .A1(n5933), .A2(n5872), .B1(n5933), .B2(SRAM_out_buffer[44]), 
        .O(n3114) );
  MOAI1S U6768 ( .A1(n5934), .A2(n5872), .B1(n5934), .B2(SRAM_out_buffer[76]), 
        .O(n3113) );
  MOAI1S U6769 ( .A1(n5934), .A2(n5878), .B1(n5934), .B2(SRAM_out_buffer[78]), 
        .O(n3101) );
  MOAI1S U6770 ( .A1(n5934), .A2(n5857), .B1(n5934), .B2(SRAM_out_buffer[79]), 
        .O(n3095) );
  FA1S U6771 ( .A(n5861), .B(n5864), .CI(pool_temp[17]), .CO(n5774) );
  ND2S U6772 ( .I1(pool_temp[23]), .I2(n5780), .O(n5779) );
  MOAI1S U6773 ( .A1(pool_temp[23]), .A2(n5780), .B1(n5850), .B2(n5779), .O(
        n5781) );
  INV1S U6774 ( .I(n5994), .O(n5788) );
  ND2 U6775 ( .I1(n5790), .I2(n5817), .O(n5827) );
  INV1S U6776 ( .I(pool_temp[23]), .O(n5818) );
  AOI22S U6777 ( .A1(n5875), .A2(n5791), .B1(n5878), .B2(n5813), .O(n5796) );
  AOI22S U6778 ( .A1(n5873), .A2(n5798), .B1(n5870), .B2(n5797), .O(n5803) );
  AOI22S U6779 ( .A1(n5861), .A2(n5805), .B1(n5864), .B2(n5804), .O(n5810) );
  AOI22S U6780 ( .A1(n5863), .A2(n5807), .B1(n5866), .B2(n5806), .O(n5809) );
  NR2 U6781 ( .I1(n5810), .I2(n5830), .O(n5811) );
  NR2 U6782 ( .I1(n5833), .I2(n5811), .O(n5812) );
  NR2 U6783 ( .I1(n5831), .I2(n5812), .O(n5815) );
  NR2 U6784 ( .I1(n5878), .I2(n5813), .O(n5814) );
  NR2 U6785 ( .I1(n5815), .I2(n5829), .O(n5854) );
  OAI12HS U6786 ( .B1(n5985), .B2(n5816), .A1(n5854), .O(n5826) );
  OR2 U6787 ( .I1(n5817), .I2(n5854), .O(n5825) );
  OAI222S U6788 ( .A1(n5827), .A2(n5818), .B1(n5858), .B2(n5826), .C1(n5825), 
        .C2(n5857), .O(n3092) );
  INV1S U6789 ( .I(pool_temp[16]), .O(n5819) );
  OAI222S U6790 ( .A1(n5827), .A2(n5819), .B1(n5861), .B2(n5826), .C1(n5825), 
        .C2(n5860), .O(n3090) );
  INV1S U6791 ( .I(pool_temp[17]), .O(n5820) );
  OAI222S U6792 ( .A1(n5820), .A2(n5827), .B1(n5864), .B2(n5826), .C1(n5825), 
        .C2(n5863), .O(n3088) );
  INV1S U6793 ( .I(pool_temp[18]), .O(n5821) );
  OAI222S U6794 ( .A1(n5821), .A2(n5827), .B1(n5867), .B2(n5826), .C1(n5825), 
        .C2(n5866), .O(n3086) );
  INV1S U6795 ( .I(pool_temp[19]), .O(n5822) );
  OAI222S U6796 ( .A1(n5822), .A2(n5827), .B1(n5870), .B2(n5826), .C1(n5825), 
        .C2(n5869), .O(n3084) );
  INV1S U6797 ( .I(pool_temp[20]), .O(n5823) );
  OAI222S U6798 ( .A1(n5823), .A2(n5827), .B1(n5873), .B2(n5826), .C1(n5825), 
        .C2(n5872), .O(n3082) );
  INV1S U6799 ( .I(pool_temp[21]), .O(n5824) );
  OAI222S U6800 ( .A1(n5824), .A2(n5827), .B1(n5876), .B2(n5826), .C1(n5825), 
        .C2(n5875), .O(n3080) );
  INV1S U6801 ( .I(pool_temp[22]), .O(n5828) );
  OAI222S U6802 ( .A1(n5828), .A2(n5827), .B1(n5881), .B2(n5826), .C1(n5825), 
        .C2(n5878), .O(n3078) );
  INV1S U6803 ( .I(pool_temp[7]), .O(n5859) );
  INV1S U6804 ( .I(n5829), .O(n5832) );
  MOAI1S U6805 ( .A1(n5834), .A2(n5833), .B1(n5832), .B2(n5831), .O(n5841) );
  FA1S U6806 ( .A(pool_temp[7]), .B(n5857), .CI(n5839), .CO(n5840) );
  NR2 U6807 ( .I1(n5841), .I2(n5840), .O(n5842) );
  OAI12HS U6808 ( .B1(cal_count_5[2]), .B2(n5842), .A1(n6028), .O(n5856) );
  FA1S U6809 ( .A(n5861), .B(n5864), .CI(pool_temp[1]), .CO(n5843) );
  FA1S U6810 ( .A(pool_temp[2]), .B(n5867), .CI(n5843), .CO(n5844) );
  FA1S U6811 ( .A(n5870), .B(pool_temp[3]), .CI(n5844), .CO(n5845) );
  FA1S U6812 ( .A(pool_temp[4]), .B(n5873), .CI(n5845), .CO(n5846) );
  FA1S U6813 ( .A(n5876), .B(pool_temp[5]), .CI(n5846), .CO(n5847) );
  ND2S U6814 ( .I1(pool_temp[7]), .I2(n5848), .O(n5849) );
  MOAI1S U6815 ( .A1(pool_temp[7]), .A2(n5848), .B1(n5850), .B2(n5849), .O(
        n5851) );
  ND3S U6816 ( .I1(n6028), .I2(n5854), .I3(n5851), .O(n5852) );
  INV1S U6817 ( .I(n5852), .O(n5853) );
  OAI222S U6818 ( .A1(n5859), .A2(n5882), .B1(n5858), .B2(n5880), .C1(n5879), 
        .C2(n5857), .O(n3076) );
  INV1S U6819 ( .I(pool_temp[0]), .O(n5862) );
  OAI222S U6820 ( .A1(n5882), .A2(n5862), .B1(n5861), .B2(n5880), .C1(n5879), 
        .C2(n5860), .O(n3074) );
  INV1S U6821 ( .I(pool_temp[1]), .O(n5865) );
  OAI222S U6822 ( .A1(n5865), .A2(n5882), .B1(n5864), .B2(n5880), .C1(n5879), 
        .C2(n5863), .O(n3072) );
  INV1S U6823 ( .I(pool_temp[2]), .O(n5868) );
  OAI222S U6824 ( .A1(n5868), .A2(n5882), .B1(n5867), .B2(n5880), .C1(n5879), 
        .C2(n5866), .O(n3070) );
  INV1S U6825 ( .I(pool_temp[3]), .O(n5871) );
  OAI222S U6826 ( .A1(n5871), .A2(n5882), .B1(n5870), .B2(n5880), .C1(n5879), 
        .C2(n5869), .O(n3068) );
  INV1S U6827 ( .I(pool_temp[4]), .O(n5874) );
  OAI222S U6828 ( .A1(n5874), .A2(n5882), .B1(n5873), .B2(n5880), .C1(n5879), 
        .C2(n5872), .O(n3066) );
  INV1S U6829 ( .I(pool_temp[5]), .O(n5877) );
  OAI222S U6830 ( .A1(n5877), .A2(n5882), .B1(n5876), .B2(n5880), .C1(n5879), 
        .C2(n5875), .O(n3064) );
  INV1S U6831 ( .I(pool_temp[6]), .O(n5883) );
  OAI222S U6832 ( .A1(n5883), .A2(n5882), .B1(n5881), .B2(n5880), .C1(n5879), 
        .C2(n5878), .O(n3062) );
  MOAI1S U6833 ( .A1(n5933), .A2(n6031), .B1(n5933), .B2(SRAM_out_buffer[48]), 
        .O(n3058) );
  MOAI1S U6834 ( .A1(n5934), .A2(n6031), .B1(n5934), .B2(SRAM_out_buffer[80]), 
        .O(n3057) );
  MOAI1S U6835 ( .A1(n5933), .A2(n6034), .B1(n5933), .B2(SRAM_out_buffer[49]), 
        .O(n3052) );
  MOAI1S U6836 ( .A1(n5934), .A2(n6034), .B1(n5934), .B2(SRAM_out_buffer[81]), 
        .O(n3051) );
  INV1S U6837 ( .I(n6034), .O(n5960) );
  MOAI1S U6838 ( .A1(n5934), .A2(n6037), .B1(n5934), .B2(SRAM_out_buffer[82]), 
        .O(n3045) );
  MOAI1S U6839 ( .A1(n5933), .A2(n6040), .B1(n5933), .B2(SRAM_out_buffer[51]), 
        .O(n3040) );
  MOAI1S U6840 ( .A1(n5934), .A2(n6040), .B1(n5934), .B2(SRAM_out_buffer[83]), 
        .O(n3039) );
  MOAI1S U6841 ( .A1(n5933), .A2(n6043), .B1(n5933), .B2(SRAM_out_buffer[52]), 
        .O(n3034) );
  MOAI1S U6842 ( .A1(n5934), .A2(n6043), .B1(n5934), .B2(SRAM_out_buffer[84]), 
        .O(n3033) );
  MOAI1S U6843 ( .A1(n5933), .A2(n6046), .B1(n5933), .B2(SRAM_out_buffer[53]), 
        .O(n3028) );
  MOAI1S U6844 ( .A1(n5934), .A2(n6046), .B1(n5934), .B2(SRAM_out_buffer[85]), 
        .O(n3027) );
  MOAI1S U6845 ( .A1(n5933), .A2(n6049), .B1(n5933), .B2(SRAM_out_buffer[54]), 
        .O(n3022) );
  MOAI1S U6846 ( .A1(n5934), .A2(n6049), .B1(n5934), .B2(SRAM_out_buffer[86]), 
        .O(n3021) );
  MOAI1S U6847 ( .A1(n5934), .A2(n6029), .B1(n5934), .B2(SRAM_out_buffer[87]), 
        .O(n3015) );
  MOAI1S U6848 ( .A1(n5933), .A2(n6032), .B1(n5933), .B2(SRAM_out_buffer[56]), 
        .O(n3010) );
  MOAI1S U6849 ( .A1(n5934), .A2(n6032), .B1(n5934), .B2(SRAM_out_buffer[88]), 
        .O(n3009) );
  MOAI1S U6850 ( .A1(n5933), .A2(n6035), .B1(n5933), .B2(SRAM_out_buffer[57]), 
        .O(n2998) );
  MOAI1S U6851 ( .A1(n5934), .A2(n6035), .B1(n5934), .B2(SRAM_out_buffer[89]), 
        .O(n2997) );
  OAI222S U6852 ( .A1(n6062), .A2(n5889), .B1(n6060), .B2(n6035), .C1(n5888), 
        .C2(n6057), .O(n2990) );
  INV1S U6853 ( .I(n5961), .O(n6038) );
  MOAI1S U6854 ( .A1(n5933), .A2(n6038), .B1(n5933), .B2(SRAM_out_buffer[58]), 
        .O(n2986) );
  MOAI1S U6855 ( .A1(n5934), .A2(n6038), .B1(n5934), .B2(SRAM_out_buffer[90]), 
        .O(n2985) );
  MOAI1S U6856 ( .A1(n5933), .A2(n6041), .B1(n5933), .B2(SRAM_out_buffer[59]), 
        .O(n2974) );
  MOAI1S U6857 ( .A1(n5934), .A2(n6041), .B1(n5934), .B2(SRAM_out_buffer[91]), 
        .O(n2973) );
  MOAI1S U6858 ( .A1(n5942), .A2(n5890), .B1(n5935), .B2(SRAM_out_buffer[91]), 
        .O(n5891) );
  INV1S U6859 ( .I(SRAM_out_buffer[91]), .O(n5896) );
  OAI222S U6860 ( .A1(n5893), .A2(n5943), .B1(n5896), .B2(n5941), .C1(n5895), 
        .C2(n5942), .O(n2968) );
  OAI222S U6861 ( .A1(n5896), .A2(n5946), .B1(n5895), .B2(n5943), .C1(n5894), 
        .C2(n5942), .O(n2967) );
  OAI222S U6862 ( .A1(n6062), .A2(n5898), .B1(n6060), .B2(n6041), .C1(n5897), 
        .C2(n6057), .O(n2966) );
  MOAI1S U6863 ( .A1(n5933), .A2(n6044), .B1(n5933), .B2(SRAM_out_buffer[60]), 
        .O(n2962) );
  MOAI1S U6864 ( .A1(n5934), .A2(n6044), .B1(n5934), .B2(SRAM_out_buffer[92]), 
        .O(n2961) );
  MOAI1S U6865 ( .A1(n5942), .A2(n5899), .B1(n5935), .B2(SRAM_out_buffer[92]), 
        .O(n5900) );
  OAI222S U6866 ( .A1(n5904), .A2(n5943), .B1(n5903), .B2(n5941), .C1(n5902), 
        .C2(n5942), .O(n2956) );
  OAI112HS U6867 ( .C1(n5942), .C2(n5909), .A1(n5908), .B1(n5907), .O(n2951)
         );
  MOAI1S U6868 ( .A1(n5933), .A2(n6047), .B1(n5933), .B2(SRAM_out_buffer[61]), 
        .O(n2950) );
  MOAI1S U6869 ( .A1(n5934), .A2(n6047), .B1(n5934), .B2(SRAM_out_buffer[93]), 
        .O(n2949) );
  MOAI1S U6870 ( .A1(n5942), .A2(n5910), .B1(n5935), .B2(SRAM_out_buffer[93]), 
        .O(n5911) );
  INV1S U6871 ( .I(SRAM_out_buffer[93]), .O(n5915) );
  OAI222S U6872 ( .A1(n6321), .A2(n5943), .B1(n5915), .B2(n5941), .C1(n5914), 
        .C2(n5942), .O(n2944) );
  OAI222S U6873 ( .A1(n5915), .A2(n5946), .B1(n5914), .B2(n5943), .C1(n5913), 
        .C2(n5942), .O(n2943) );
  OAI112HS U6874 ( .C1(n6068), .C2(n5922), .A1(n5921), .B1(n5920), .O(n2939)
         );
  INV1S U6875 ( .I(n5967), .O(n6052) );
  MOAI1S U6876 ( .A1(n5933), .A2(n6052), .B1(n5933), .B2(SRAM_out_buffer[62]), 
        .O(n2938) );
  MOAI1S U6877 ( .A1(n5934), .A2(n6052), .B1(n5934), .B2(SRAM_out_buffer[94]), 
        .O(n2937) );
  MOAI1S U6878 ( .A1(n5942), .A2(n5923), .B1(n5935), .B2(SRAM_out_buffer[94]), 
        .O(n5924) );
  INV1S U6879 ( .I(SRAM_out_buffer[94]), .O(n5929) );
  OAI222S U6880 ( .A1(n5928), .A2(n5942), .B1(n5929), .B2(n5941), .C1(n5926), 
        .C2(n5943), .O(n2932) );
  OAI222S U6881 ( .A1(n5929), .A2(n5946), .B1(n5928), .B2(n5943), .C1(n5927), 
        .C2(n5942), .O(n2931) );
  MOAI1S U6882 ( .A1(n5933), .A2(n6059), .B1(n5933), .B2(SRAM_out_buffer[63]), 
        .O(n2926) );
  MOAI1S U6883 ( .A1(n5934), .A2(n6059), .B1(n5934), .B2(SRAM_out_buffer[95]), 
        .O(n2925) );
  MOAI1S U6884 ( .A1(n5942), .A2(n5936), .B1(n5935), .B2(SRAM_out_buffer[95]), 
        .O(n5937) );
  INV1S U6885 ( .I(SRAM_out_buffer[95]), .O(n5947) );
  OAI222S U6886 ( .A1(n5944), .A2(n5942), .B1(n5947), .B2(n5941), .C1(n5940), 
        .C2(n5943), .O(n2920) );
  OAI222S U6887 ( .A1(n5947), .A2(n5946), .B1(n5945), .B2(n5942), .C1(n5944), 
        .C2(n5943), .O(n2919) );
  AOI22S U6888 ( .A1(n6052), .A2(n5949), .B1(n6047), .B2(n5948), .O(n5954) );
  AOI22S U6889 ( .A1(n6040), .A2(n5956), .B1(n6043), .B2(n5955), .O(n5959) );
  NR2 U6890 ( .I1(n5956), .I2(n6040), .O(n5963) );
  OR3B2S U6891 ( .I1(n5963), .B1(n6037), .B2(n5961), .O(n5957) );
  MOAI1S U6892 ( .A1(n6037), .A2(n5961), .B1(n6035), .B2(n5960), .O(n5962) );
  NR2 U6893 ( .I1(n5963), .I2(n5962), .O(n5971) );
  MOAI1S U6894 ( .A1(n5965), .A2(n6035), .B1(n5971), .B2(n5964), .O(n5966) );
  NR2 U6895 ( .I1(n5972), .I2(n5966), .O(n5970) );
  INV1S U6896 ( .I(n6027), .O(n6014) );
  NR2 U6897 ( .I1(n5972), .I2(n5971), .O(n5975) );
  FA1S U6898 ( .A(n6032), .B(n6035), .CI(pool_temp[25]), .CO(n5976) );
  NR2 U6899 ( .I1(n6013), .I2(n5982), .O(n5983) );
  AOI22H U6900 ( .A1(n5985), .A2(n6014), .B1(n5984), .B2(n5983), .O(n6003) );
  FA1S U6901 ( .A(pool_temp[25]), .B(n6034), .CI(n6031), .CO(n5986) );
  FA1S U6902 ( .A(n6037), .B(pool_temp[26]), .CI(n5986), .CO(n5987) );
  FA1S U6903 ( .A(pool_temp[27]), .B(n6040), .CI(n5987), .CO(n5988) );
  FA1S U6904 ( .A(pool_temp[28]), .B(n6043), .CI(n5988), .CO(n5989) );
  FA1S U6905 ( .A(pool_temp[29]), .B(n6046), .CI(n5989), .CO(n5990) );
  ND2S U6906 ( .I1(n5992), .I2(cal_count_5[0]), .O(n5993) );
  ND3P U6907 ( .I1(n6027), .I2(n5994), .I3(n5993), .O(n6002) );
  INV1S U6908 ( .I(pool_temp[31]), .O(n5995) );
  OAI222S U6909 ( .A1(n6004), .A2(n5995), .B1(n6059), .B2(n6003), .C1(n6002), 
        .C2(n6029), .O(n2918) );
  INV1S U6910 ( .I(pool_temp[24]), .O(n5996) );
  OAI222S U6911 ( .A1(n6004), .A2(n5996), .B1(n6032), .B2(n6003), .C1(n6002), 
        .C2(n6031), .O(n2917) );
  INV1S U6912 ( .I(pool_temp[25]), .O(n5997) );
  OAI222S U6913 ( .A1(n5997), .A2(n6004), .B1(n6035), .B2(n6003), .C1(n6002), 
        .C2(n6034), .O(n2915) );
  INV1S U6914 ( .I(pool_temp[26]), .O(n5998) );
  OAI222S U6915 ( .A1(n5998), .A2(n6004), .B1(n6038), .B2(n6003), .C1(n6002), 
        .C2(n6037), .O(n2913) );
  INV1S U6916 ( .I(pool_temp[27]), .O(n5999) );
  OAI222S U6917 ( .A1(n5999), .A2(n6004), .B1(n6041), .B2(n6003), .C1(n6002), 
        .C2(n6040), .O(n2911) );
  INV1S U6918 ( .I(pool_temp[28]), .O(n6000) );
  OAI222S U6919 ( .A1(n6000), .A2(n6004), .B1(n6044), .B2(n6003), .C1(n6002), 
        .C2(n6043), .O(n2909) );
  INV1S U6920 ( .I(pool_temp[29]), .O(n6001) );
  OAI222S U6921 ( .A1(n6001), .A2(n6004), .B1(n6047), .B2(n6003), .C1(n6002), 
        .C2(n6046), .O(n2907) );
  INV1S U6922 ( .I(pool_temp[30]), .O(n6005) );
  OAI222S U6923 ( .A1(n6005), .A2(n6004), .B1(n6052), .B2(n6003), .C1(n6002), 
        .C2(n6049), .O(n2905) );
  INV1S U6924 ( .I(pool_temp[15]), .O(n6030) );
  FA1S U6925 ( .A(n6032), .B(n6035), .CI(pool_temp[9]), .CO(n6006) );
  NR2 U6926 ( .I1(n6013), .I2(n6012), .O(n6017) );
  FA1S U6927 ( .A(pool_temp[9]), .B(n6034), .CI(pool_temp[8]), .CO(n6018) );
  ND2S U6928 ( .I1(n6025), .I2(n6024), .O(n6026) );
  OAI222S U6929 ( .A1(n6030), .A2(n6053), .B1(n6059), .B2(n6051), .C1(n6050), 
        .C2(n6029), .O(n2903) );
  INV1S U6930 ( .I(pool_temp[8]), .O(n6033) );
  OAI222S U6931 ( .A1(n6033), .A2(n6053), .B1(n6032), .B2(n6051), .C1(n6050), 
        .C2(n6031), .O(n2901) );
  INV1S U6932 ( .I(pool_temp[9]), .O(n6036) );
  OAI222S U6933 ( .A1(n6036), .A2(n6053), .B1(n6035), .B2(n6051), .C1(n6050), 
        .C2(n6034), .O(n2899) );
  INV1S U6934 ( .I(pool_temp[10]), .O(n6039) );
  OAI222S U6935 ( .A1(n6039), .A2(n6053), .B1(n6038), .B2(n6051), .C1(n6050), 
        .C2(n6037), .O(n2897) );
  INV1S U6936 ( .I(pool_temp[11]), .O(n6042) );
  OAI222S U6937 ( .A1(n6042), .A2(n6053), .B1(n6041), .B2(n6051), .C1(n6050), 
        .C2(n6040), .O(n2895) );
  INV1S U6938 ( .I(pool_temp[12]), .O(n6045) );
  OAI222S U6939 ( .A1(n6045), .A2(n6053), .B1(n6044), .B2(n6051), .C1(n6050), 
        .C2(n6043), .O(n2893) );
  INV1S U6940 ( .I(pool_temp[13]), .O(n6048) );
  OAI222S U6941 ( .A1(n6048), .A2(n6053), .B1(n6047), .B2(n6051), .C1(n6050), 
        .C2(n6046), .O(n2891) );
  INV1S U6942 ( .I(pool_temp[14]), .O(n6054) );
  OAI222S U6943 ( .A1(n6054), .A2(n6053), .B1(n6052), .B2(n6051), .C1(n6050), 
        .C2(n6049), .O(n2889) );
  OAI222S U6944 ( .A1(n6062), .A2(n6061), .B1(n6060), .B2(n6059), .C1(n6058), 
        .C2(n6057), .O(n2887) );
  AOI22S U6945 ( .A1(median_in[23]), .A2(n6064), .B1(n3517), .B2(n6063), .O(
        n6066) );
  OAI112HS U6946 ( .C1(n6068), .C2(n6067), .A1(n6066), .B1(n6065), .O(n2884)
         );
  ND2S U6947 ( .I1(n6069), .I2(conv_out_reg[16]), .O(n6076) );
  ND3S U6948 ( .I1(wait_conv_out_count[1]), .I2(conv_out_reg[17]), .I3(n6302), 
        .O(n6075) );
  ND3S U6949 ( .I1(n6070), .I2(wait_conv_out_count[0]), .I3(conv_out_reg[18]), 
        .O(n6074) );
  INV1S U6950 ( .I(conv_out_reg[19]), .O(n6072) );
  NR2 U6951 ( .I1(n6072), .I2(n6071), .O(n6073) );
  AN4B1S U6952 ( .I1(n6076), .I2(n6075), .I3(n6074), .B1(n6073), .O(n61180) );
  AOI22S U6953 ( .A1(n6094), .A2(conv_out_reg[2]), .B1(n6093), .B2(
        conv_out_reg[0]), .O(n6078) );
  ND2S U6954 ( .I1(n6090), .I2(conv_out_reg[4]), .O(n6077) );
  ND3S U6955 ( .I1(n6078), .I2(wait_conv_out_count[0]), .I3(n6077), .O(n6104)
         );
  ND2S U6956 ( .I1(n6093), .I2(conv_out_reg[1]), .O(n6103) );
  INV1S U6957 ( .I(conv_out_reg[7]), .O(n6079) );
  ND2S U6958 ( .I1(n6103), .I2(n6079), .O(n6082) );
  ND2S U6959 ( .I1(n6090), .I2(conv_out_reg[5]), .O(n6081) );
  ND2S U6960 ( .I1(n6094), .I2(conv_out_reg[3]), .O(n6080) );
  ND3S U6961 ( .I1(n6081), .I2(n6302), .I3(n6080), .O(n6106) );
  OAI22S U6962 ( .A1(conv_out_reg[6]), .A2(n6104), .B1(n6082), .B2(n6106), .O(
        n6085) );
  ND2S U6963 ( .I1(n6084), .I2(n6083), .O(n6109) );
  ND2S U6964 ( .I1(n6085), .I2(n6109), .O(n6113) );
  INV1S U6965 ( .I(n6090), .O(n6087) );
  INV1S U6966 ( .I(conv_out_reg[12]), .O(n6086) );
  MOAI1S U6967 ( .A1(n6087), .A2(n6086), .B1(n6093), .B2(conv_out_reg[8]), .O(
        n6100) );
  ND2S U6968 ( .I1(n6107), .I2(conv_out_reg[14]), .O(n6089) );
  ND2S U6969 ( .I1(n6094), .I2(conv_out_reg[10]), .O(n6088) );
  ND2S U6970 ( .I1(n6090), .I2(conv_out_reg[13]), .O(n6092) );
  ND2S U6971 ( .I1(n6107), .I2(conv_out_reg[15]), .O(n6091) );
  ND3S U6972 ( .I1(n6092), .I2(n6302), .I3(n6091), .O(n6098) );
  INV1S U6973 ( .I(n6093), .O(n6096) );
  INV1S U6974 ( .I(conv_out_reg[9]), .O(n6095) );
  MOAI1S U6975 ( .A1(n6096), .A2(n6095), .B1(n6094), .B2(conv_out_reg[11]), 
        .O(n6097) );
  OAI22S U6976 ( .A1(n6100), .A2(n6099), .B1(n6098), .B2(n6097), .O(n6102) );
  INV1S U6977 ( .I(n6109), .O(n6101) );
  ND2S U6978 ( .I1(n6102), .I2(n6101), .O(n6112) );
  INV1S U6979 ( .I(n6103), .O(n6105) );
  OAI12HS U6980 ( .B1(n6106), .B2(n6105), .A1(n6104), .O(n6110) );
  INV1S U6981 ( .I(n6107), .O(n6108) );
  ND3S U6982 ( .I1(n6113), .I2(n6112), .I3(n6111), .O(n61170) );
  OAI12HS U6983 ( .B1(wait_conv_out_count[4]), .B2(n61150), .A1(n6114), .O(
        n61160) );
  MUX2S U6984 ( .A(n61180), .B(n61170), .S(n61160), .O(n61210) );
  INV1S U6985 ( .I(out_value), .O(n61200) );
  MUX2S U6986 ( .A(n61210), .B(n61200), .S(n61190), .O(n61220) );
  NR2 U6987 ( .I1(n61230), .I2(n61220), .O(n2864) );
  INV1S U6988 ( .I(n61240), .O(n61270) );
  MOAI1S U6989 ( .A1(n61270), .A2(n61250), .B1(n61270), .B2(image_size[0]), 
        .O(n2861) );
  MOAI1S U6990 ( .A1(n61270), .A2(n61260), .B1(n61270), .B2(image_size[1]), 
        .O(n2860) );
  MOAI1S U6991 ( .A1(n3491), .A2(n61280), .B1(n3491), .B2(conv_out_reg[0]), 
        .O(n2859) );
  MOAI1S U6992 ( .A1(n3491), .A2(n61290), .B1(n3491), .B2(conv_out_reg[17]), 
        .O(n2856) );
  MOAI1S U6993 ( .A1(n3491), .A2(n61300), .B1(n3491), .B2(conv_out_reg[16]), 
        .O(n2855) );
  MOAI1S U6994 ( .A1(n3491), .A2(n6131), .B1(n3491), .B2(conv_out_reg[15]), 
        .O(n2854) );
  MOAI1S U6995 ( .A1(n3491), .A2(n6132), .B1(n3491), .B2(conv_out_reg[14]), 
        .O(n2853) );
  MOAI1S U6996 ( .A1(n3491), .A2(n6133), .B1(n3491), .B2(conv_out_reg[13]), 
        .O(n2852) );
  MOAI1S U6997 ( .A1(n3491), .A2(n6134), .B1(n3491), .B2(conv_out_reg[12]), 
        .O(n2851) );
  MOAI1S U6998 ( .A1(n3491), .A2(n6135), .B1(n3491), .B2(conv_out_reg[11]), 
        .O(n2850) );
  MOAI1S U6999 ( .A1(n3491), .A2(n6136), .B1(n3491), .B2(conv_out_reg[10]), 
        .O(n2849) );
  MOAI1S U7000 ( .A1(n3491), .A2(n6137), .B1(n3491), .B2(conv_out_reg[9]), .O(
        n2848) );
  MOAI1S U7001 ( .A1(n3491), .A2(n6138), .B1(n3491), .B2(conv_out_reg[8]), .O(
        n2847) );
  MOAI1S U7002 ( .A1(n3491), .A2(n6139), .B1(n3491), .B2(conv_out_reg[7]), .O(
        n2846) );
  MOAI1S U7003 ( .A1(n3491), .A2(n6140), .B1(n3491), .B2(conv_out_reg[6]), .O(
        n2845) );
  MOAI1S U7004 ( .A1(n3491), .A2(n6141), .B1(n3491), .B2(conv_out_reg[5]), .O(
        n2844) );
  MOAI1S U7005 ( .A1(n3491), .A2(n6142), .B1(n3491), .B2(conv_out_reg[4]), .O(
        n2843) );
  MOAI1S U7006 ( .A1(n3491), .A2(n6143), .B1(n3491), .B2(conv_out_reg[3]), .O(
        n2842) );
  MOAI1S U7007 ( .A1(n3491), .A2(n3504), .B1(n3491), .B2(conv_out_reg[2]), .O(
        n2841) );
  MOAI1S U7008 ( .A1(n3491), .A2(n6144), .B1(n3491), .B2(conv_out_reg[1]), .O(
        n2840) );
  INV1S U7009 ( .I(gray_wgt_reg[31]), .O(n6160) );
  MAOI1S U7010 ( .A1(n6145), .A2(wgt_temp[7]), .B1(n6145), .B2(wgt_temp[7]), 
        .O(n6146) );
  INV1S U7011 ( .I(gray_wgt_reg[30]), .O(n6161) );
  HA1 U7012 ( .A(wgt_temp[6]), .B(n6147), .C(n6145), .S(n6148) );
  MOAI1S U7013 ( .A1(n6196), .A2(n6161), .B1(n6196), .B2(n6148), .O(n2838) );
  INV1S U7014 ( .I(gray_wgt_reg[29]), .O(n6162) );
  FA1S U7015 ( .A(image[7]), .B(wgt_temp[5]), .CI(n6149), .CO(n6147), .S(n6150) );
  MOAI1S U7016 ( .A1(n6196), .A2(n6162), .B1(n6196), .B2(n6150), .O(n2837) );
  INV1S U7017 ( .I(gray_wgt_reg[28]), .O(n6163) );
  FA1S U7018 ( .A(image[6]), .B(wgt_temp[4]), .CI(n6151), .CO(n6149), .S(n6152) );
  MOAI1S U7019 ( .A1(n6196), .A2(n6163), .B1(n6196), .B2(n6152), .O(n2836) );
  INV1S U7020 ( .I(gray_wgt_reg[27]), .O(n6164) );
  FA1S U7021 ( .A(image[5]), .B(wgt_temp[3]), .CI(n6153), .CO(n6151), .S(n6154) );
  MOAI1S U7022 ( .A1(n6196), .A2(n6164), .B1(n6196), .B2(n6154), .O(n2835) );
  INV1S U7023 ( .I(gray_wgt_reg[26]), .O(n6165) );
  FA1S U7024 ( .A(image[4]), .B(wgt_temp[2]), .CI(n6155), .CO(n6153), .S(n6156) );
  MOAI1S U7025 ( .A1(n6196), .A2(n6165), .B1(n6196), .B2(n6156), .O(n2834) );
  INV1S U7026 ( .I(gray_wgt_reg[25]), .O(n6166) );
  FA1S U7027 ( .A(image[3]), .B(wgt_temp[1]), .CI(n6157), .CO(n6155), .S(n6158) );
  MOAI1S U7028 ( .A1(n6196), .A2(n6166), .B1(n6196), .B2(n6158), .O(n2833) );
  INV1S U7029 ( .I(gray_wgt_reg[24]), .O(n6167) );
  MOAI1S U7030 ( .A1(n6196), .A2(n6167), .B1(n6196), .B2(n6159), .O(n2832) );
  MOAI1S U7031 ( .A1(n6177), .A2(n6160), .B1(n6188), .B2(gray_wgt_reg[23]), 
        .O(n2831) );
  MOAI1S U7032 ( .A1(n6177), .A2(n6161), .B1(n6193), .B2(gray_wgt_reg[22]), 
        .O(n2830) );
  INV1S U7033 ( .I(n6196), .O(n6188) );
  INV1S U7034 ( .I(n6196), .O(n6193) );
  MOAI1S U7035 ( .A1(n6188), .A2(n6162), .B1(n6193), .B2(gray_wgt_reg[21]), 
        .O(n2829) );
  MOAI1S U7036 ( .A1(n6188), .A2(n6163), .B1(n6193), .B2(gray_wgt_reg[20]), 
        .O(n2828) );
  MOAI1S U7037 ( .A1(n6177), .A2(n6164), .B1(n6193), .B2(gray_wgt_reg[19]), 
        .O(n2827) );
  MOAI1S U7038 ( .A1(n6188), .A2(n6165), .B1(n6193), .B2(gray_wgt_reg[18]), 
        .O(n2826) );
  INV1S U7039 ( .I(n6196), .O(n6177) );
  MOAI1S U7040 ( .A1(n6193), .A2(n6166), .B1(n6177), .B2(gray_wgt_reg[17]), 
        .O(n2825) );
  MOAI1S U7041 ( .A1(n6193), .A2(n6167), .B1(n6177), .B2(gray_wgt_reg[16]), 
        .O(n2824) );
  INV1S U7042 ( .I(gray_wgt_reg[15]), .O(n6169) );
  MOAI1S U7043 ( .A1(n6196), .A2(n6169), .B1(n6196), .B2(gray_wgt_reg[23]), 
        .O(n2823) );
  INV1S U7044 ( .I(gray_wgt_reg[14]), .O(n6170) );
  MOAI1S U7045 ( .A1(n6196), .A2(n6170), .B1(n6196), .B2(gray_wgt_reg[22]), 
        .O(n2822) );
  INV1S U7046 ( .I(gray_wgt_reg[13]), .O(n6171) );
  MOAI1S U7047 ( .A1(n6196), .A2(n6171), .B1(n6196), .B2(gray_wgt_reg[21]), 
        .O(n2821) );
  INV1S U7048 ( .I(gray_wgt_reg[12]), .O(n6172) );
  MOAI1S U7049 ( .A1(n6196), .A2(n6172), .B1(n6196), .B2(gray_wgt_reg[20]), 
        .O(n2820) );
  INV1S U7050 ( .I(gray_wgt_reg[11]), .O(n6173) );
  MOAI1S U7051 ( .A1(n6196), .A2(n6173), .B1(n6196), .B2(gray_wgt_reg[19]), 
        .O(n2819) );
  INV1S U7052 ( .I(gray_wgt_reg[10]), .O(n6174) );
  MOAI1S U7053 ( .A1(n6196), .A2(n6174), .B1(n6196), .B2(gray_wgt_reg[18]), 
        .O(n2818) );
  INV1S U7054 ( .I(gray_wgt_reg[9]), .O(n6175) );
  MOAI1S U7055 ( .A1(n6196), .A2(n6175), .B1(n6196), .B2(gray_wgt_reg[17]), 
        .O(n2817) );
  INV1S U7056 ( .I(gray_wgt_reg[8]), .O(n6168) );
  MOAI1S U7057 ( .A1(n6196), .A2(n6168), .B1(n6196), .B2(gray_wgt_reg[16]), 
        .O(n2816) );
  MOAI1S U7058 ( .A1(n6193), .A2(n6168), .B1(n6177), .B2(gray_wgt_reg[0]), .O(
        n2815) );
  MOAI1S U7059 ( .A1(n6188), .A2(n6169), .B1(n6177), .B2(gray_wgt_reg[7]), .O(
        n2814) );
  MOAI1S U7060 ( .A1(n6188), .A2(n6170), .B1(n6177), .B2(gray_wgt_reg[6]), .O(
        n2813) );
  MOAI1S U7061 ( .A1(n6177), .A2(n6171), .B1(n6177), .B2(gray_wgt_reg[5]), .O(
        n2812) );
  MOAI1S U7062 ( .A1(n6188), .A2(n6172), .B1(n6177), .B2(gray_wgt_reg[4]), .O(
        n2811) );
  MOAI1S U7063 ( .A1(n6193), .A2(n6173), .B1(n6177), .B2(gray_wgt_reg[3]), .O(
        n2810) );
  MOAI1S U7064 ( .A1(n6188), .A2(n6174), .B1(n6177), .B2(gray_wgt_reg[2]), .O(
        n2809) );
  MOAI1S U7065 ( .A1(n6188), .A2(n6175), .B1(n6177), .B2(gray_wgt_reg[1]), .O(
        n2808) );
  INV1S U7066 ( .I(n6190), .O(n6191) );
  OAI22S U7067 ( .A1(n6191), .A2(max_temp[6]), .B1(n6190), .B2(image[6]), .O(
        n6176) );
  MOAI1S U7068 ( .A1(n6188), .A2(n6176), .B1(n6177), .B2(gray_max_temp[30]), 
        .O(n2807) );
  INV1S U7069 ( .I(gray_max_temp[14]), .O(n6178) );
  MOAI1S U7070 ( .A1(n6196), .A2(n6178), .B1(n6196), .B2(gray_max_temp[22]), 
        .O(n2805) );
  MOAI1S U7071 ( .A1(n6188), .A2(n6178), .B1(n6177), .B2(gray_max_temp[6]), 
        .O(n2804) );
  OAI22S U7072 ( .A1(n6191), .A2(max_temp[0]), .B1(n6190), .B2(image[0]), .O(
        n6179) );
  MOAI1S U7073 ( .A1(n6188), .A2(n6179), .B1(n6193), .B2(gray_max_temp[24]), 
        .O(n2803) );
  INV1S U7074 ( .I(gray_max_temp[8]), .O(n6180) );
  MOAI1S U7075 ( .A1(n6196), .A2(n6180), .B1(n6196), .B2(gray_max_temp[16]), 
        .O(n2801) );
  MOAI1S U7076 ( .A1(n6193), .A2(n6180), .B1(n6188), .B2(gray_max_temp[0]), 
        .O(n2800) );
  OAI22S U7077 ( .A1(n6191), .A2(max_temp[1]), .B1(n6190), .B2(image[1]), .O(
        n6181) );
  MOAI1S U7078 ( .A1(n6193), .A2(n6181), .B1(n6177), .B2(gray_max_temp[25]), 
        .O(n2799) );
  INV1S U7079 ( .I(gray_max_temp[9]), .O(n6182) );
  MOAI1S U7080 ( .A1(n6196), .A2(n6182), .B1(n6196), .B2(gray_max_temp[17]), 
        .O(n2797) );
  MOAI1S U7081 ( .A1(n6193), .A2(n6182), .B1(n6177), .B2(gray_max_temp[1]), 
        .O(n2796) );
  OAI22S U7082 ( .A1(n6191), .A2(max_temp[2]), .B1(n6190), .B2(image[2]), .O(
        n6183) );
  MOAI1S U7083 ( .A1(n6193), .A2(n6183), .B1(n6193), .B2(gray_max_temp[26]), 
        .O(n2795) );
  INV1S U7084 ( .I(gray_max_temp[10]), .O(n6184) );
  MOAI1S U7085 ( .A1(n6196), .A2(n6184), .B1(n6196), .B2(gray_max_temp[18]), 
        .O(n2793) );
  MOAI1S U7086 ( .A1(n6193), .A2(n6184), .B1(n6188), .B2(gray_max_temp[2]), 
        .O(n2792) );
  OAI22S U7087 ( .A1(n6191), .A2(max_temp[3]), .B1(n6190), .B2(image[3]), .O(
        n6185) );
  MOAI1S U7088 ( .A1(n6193), .A2(n6185), .B1(n6188), .B2(gray_max_temp[27]), 
        .O(n2791) );
  INV1S U7089 ( .I(gray_max_temp[11]), .O(n6186) );
  MOAI1S U7090 ( .A1(n6196), .A2(n6186), .B1(n6196), .B2(gray_max_temp[19]), 
        .O(n2789) );
  MOAI1S U7091 ( .A1(n6188), .A2(n6186), .B1(n6177), .B2(gray_max_temp[3]), 
        .O(n2788) );
  OAI22S U7092 ( .A1(n6191), .A2(max_temp[4]), .B1(n6190), .B2(image[4]), .O(
        n6187) );
  MOAI1S U7093 ( .A1(n6188), .A2(n6187), .B1(n6188), .B2(gray_max_temp[28]), 
        .O(n2787) );
  INV1S U7094 ( .I(gray_max_temp[12]), .O(n6189) );
  MOAI1S U7095 ( .A1(n6196), .A2(n6189), .B1(n6196), .B2(gray_max_temp[20]), 
        .O(n2785) );
  MOAI1S U7096 ( .A1(n6177), .A2(n6189), .B1(n6177), .B2(gray_max_temp[4]), 
        .O(n2784) );
  OAI22S U7097 ( .A1(n6191), .A2(max_temp[5]), .B1(n6190), .B2(image[5]), .O(
        n6192) );
  MOAI1S U7098 ( .A1(n6193), .A2(n6192), .B1(n6193), .B2(gray_max_temp[29]), 
        .O(n2783) );
  INV1S U7099 ( .I(gray_max_temp[13]), .O(n6194) );
  MOAI1S U7100 ( .A1(n6196), .A2(n6194), .B1(n6196), .B2(gray_max_temp[21]), 
        .O(n2781) );
  MOAI1S U7101 ( .A1(n6188), .A2(n6194), .B1(n6193), .B2(gray_max_temp[5]), 
        .O(n2780) );
  NR2 U7102 ( .I1(max_temp[7]), .I2(image[7]), .O(n6195) );
  MOAI1S U7103 ( .A1(n6193), .A2(n6195), .B1(n6188), .B2(gray_max_temp[31]), 
        .O(n2779) );
  INV1S U7104 ( .I(gray_max_temp[15]), .O(n6197) );
  MOAI1S U7105 ( .A1(n6196), .A2(n6197), .B1(n6196), .B2(gray_max_temp[23]), 
        .O(n2777) );
  MOAI1S U7106 ( .A1(n6188), .A2(n6197), .B1(n6177), .B2(gray_max_temp[7]), 
        .O(n2776) );
  NR2 U7107 ( .I1(avg_temp[7]), .I2(n6198), .O(n6201) );
  MOAI1S U7108 ( .A1(n6201), .A2(n6200), .B1(gray_avg_reg[31]), .B2(n6219), 
        .O(n2775) );
  INV1S U7109 ( .I(gray_avg_reg[29]), .O(n6209) );
  MOAI1S U7110 ( .A1(n6210), .A2(n6209), .B1(n6210), .B2(n6202), .O(n2773) );
  MOAI1S U7111 ( .A1(n6219), .A2(n6205), .B1(n6219), .B2(gray_avg_reg[26]), 
        .O(n2770) );
  MOAI1S U7112 ( .A1(n6219), .A2(n6209), .B1(n6219), .B2(gray_avg_reg[21]), 
        .O(n2765) );
  INV1S U7113 ( .I(gray_avg_reg[15]), .O(n6212) );
  MOAI1S U7114 ( .A1(n6210), .A2(n6212), .B1(n6210), .B2(gray_avg_reg[23]), 
        .O(n2759) );
  INV1S U7115 ( .I(gray_avg_reg[14]), .O(n6213) );
  MOAI1S U7116 ( .A1(n6210), .A2(n6213), .B1(n6210), .B2(gray_avg_reg[22]), 
        .O(n2758) );
  INV1S U7117 ( .I(gray_avg_reg[13]), .O(n6214) );
  MOAI1S U7118 ( .A1(n6210), .A2(n6214), .B1(n6210), .B2(gray_avg_reg[21]), 
        .O(n2757) );
  INV1S U7119 ( .I(gray_avg_reg[12]), .O(n6215) );
  MOAI1S U7120 ( .A1(n6210), .A2(n6215), .B1(n6210), .B2(gray_avg_reg[20]), 
        .O(n2756) );
  INV1S U7121 ( .I(gray_avg_reg[11]), .O(n6216) );
  MOAI1S U7122 ( .A1(n6210), .A2(n6216), .B1(n6210), .B2(gray_avg_reg[19]), 
        .O(n2755) );
  INV1S U7123 ( .I(gray_avg_reg[10]), .O(n6217) );
  MOAI1S U7124 ( .A1(n6210), .A2(n6217), .B1(n6210), .B2(gray_avg_reg[18]), 
        .O(n2754) );
  INV1S U7125 ( .I(gray_avg_reg[9]), .O(n6218) );
  MOAI1S U7126 ( .A1(n6210), .A2(n6218), .B1(n6210), .B2(gray_avg_reg[17]), 
        .O(n2753) );
  INV1S U7127 ( .I(gray_avg_reg[8]), .O(n6211) );
  MOAI1S U7128 ( .A1(n6210), .A2(n6211), .B1(n6210), .B2(gray_avg_reg[16]), 
        .O(n2752) );
  MOAI1S U7129 ( .A1(n6219), .A2(n6211), .B1(n6219), .B2(gray_avg_reg[0]), .O(
        n2751) );
  MOAI1S U7130 ( .A1(n6219), .A2(n6212), .B1(n6219), .B2(gray_avg_reg[7]), .O(
        n2750) );
  MOAI1S U7131 ( .A1(n6219), .A2(n6213), .B1(n6219), .B2(gray_avg_reg[6]), .O(
        n2749) );
  MOAI1S U7132 ( .A1(n6219), .A2(n6214), .B1(n6219), .B2(gray_avg_reg[5]), .O(
        n2748) );
  MOAI1S U7133 ( .A1(n6219), .A2(n6215), .B1(n6219), .B2(gray_avg_reg[4]), .O(
        n2747) );
  MOAI1S U7134 ( .A1(n6219), .A2(n6216), .B1(n6219), .B2(gray_avg_reg[3]), .O(
        n2746) );
  MOAI1S U7135 ( .A1(n6219), .A2(n6217), .B1(n6219), .B2(gray_avg_reg[2]), .O(
        n2745) );
  MOAI1S U7136 ( .A1(n6219), .A2(n6218), .B1(n6219), .B2(gray_avg_reg[1]), .O(
        n2744) );
  INV1S U7137 ( .I(SRAM_192X32_out_decode[9]), .O(n6220) );
  MOAI1S U7138 ( .A1(n6265), .A2(n6220), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_192X32_data_out[9]), .O(n2743) );
  INV1S U7139 ( .I(SRAM_192X32_out_decode[8]), .O(n6221) );
  MOAI1S U7140 ( .A1(n6265), .A2(n6221), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_192X32_data_out[8]), .O(n2742) );
  INV1S U7141 ( .I(SRAM_192X32_out_decode[7]), .O(n6222) );
  MOAI1S U7142 ( .A1(n6265), .A2(n6222), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_192X32_data_out[7]), .O(n2741) );
  INV1S U7143 ( .I(SRAM_192X32_out_decode[5]), .O(n6223) );
  MOAI1S U7144 ( .A1(n6265), .A2(n6223), .B1(n6265), .B2(
        SRAM_192X32_data_out[5]), .O(n2739) );
  INV1S U7145 ( .I(SRAM_192X32_out_decode[4]), .O(n6224) );
  MOAI1S U7146 ( .A1(n6265), .A2(n6224), .B1(n6265), .B2(
        SRAM_192X32_data_out[4]), .O(n2738) );
  INV1S U7147 ( .I(SRAM_192X32_out_decode[31]), .O(n6225) );
  MOAI1S U7148 ( .A1(n6265), .A2(n6225), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_192X32_data_out[31]), .O(n2737) );
  INV1S U7149 ( .I(SRAM_192X32_out_decode[30]), .O(n6226) );
  MOAI1S U7150 ( .A1(n6265), .A2(n6226), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_192X32_data_out[30]), .O(n2736) );
  INV1S U7151 ( .I(SRAM_192X32_out_decode[3]), .O(n6227) );
  MOAI1S U7152 ( .A1(n6265), .A2(n6227), .B1(n6265), .B2(
        SRAM_192X32_data_out[3]), .O(n2735) );
  INV1S U7153 ( .I(SRAM_192X32_out_decode[27]), .O(n6228) );
  MOAI1S U7154 ( .A1(n6265), .A2(n6228), .B1(n6265), .B2(
        SRAM_192X32_data_out[27]), .O(n2732) );
  INV1S U7155 ( .I(SRAM_192X32_out_decode[26]), .O(n6229) );
  MOAI1S U7156 ( .A1(n6265), .A2(n6229), .B1(n6265), .B2(
        SRAM_192X32_data_out[26]), .O(n2731) );
  INV1S U7157 ( .I(SRAM_192X32_out_decode[24]), .O(n6230) );
  MOAI1S U7158 ( .A1(n6265), .A2(n6230), .B1(n6265), .B2(
        SRAM_192X32_data_out[24]), .O(n2729) );
  INV1S U7159 ( .I(SRAM_192X32_out_decode[23]), .O(n6231) );
  MOAI1S U7160 ( .A1(n6265), .A2(n6231), .B1(n6265), .B2(
        SRAM_192X32_data_out[23]), .O(n2728) );
  INV1S U7161 ( .I(SRAM_192X32_out_decode[15]), .O(n6232) );
  MOAI1S U7162 ( .A1(conv_sram_stop_flag_reg), .A2(n6232), .B1(n6265), .B2(
        SRAM_192X32_data_out[15]), .O(n2719) );
  INV1S U7163 ( .I(SRAM_192X32_out_decode[14]), .O(n6233) );
  MOAI1S U7164 ( .A1(conv_sram_stop_flag_reg), .A2(n6233), .B1(n6265), .B2(
        SRAM_192X32_data_out[14]), .O(n2718) );
  INV1S U7165 ( .I(SRAM_192X32_out_decode[13]), .O(n6234) );
  MOAI1S U7166 ( .A1(conv_sram_stop_flag_reg), .A2(n6234), .B1(n6265), .B2(
        SRAM_192X32_data_out[13]), .O(n2717) );
  INV1S U7167 ( .I(SRAM_192X32_out_decode[12]), .O(n6235) );
  MOAI1S U7168 ( .A1(conv_sram_stop_flag_reg), .A2(n6235), .B1(n6265), .B2(
        SRAM_192X32_data_out[12]), .O(n2716) );
  INV1S U7169 ( .I(SRAM_192X32_out_decode[11]), .O(n6236) );
  MOAI1S U7170 ( .A1(conv_sram_stop_flag_reg), .A2(n6236), .B1(n6265), .B2(
        SRAM_192X32_data_out[11]), .O(n2715) );
  INV1S U7171 ( .I(SRAM_192X32_out_decode[10]), .O(n6237) );
  MOAI1S U7172 ( .A1(conv_sram_stop_flag_reg), .A2(n6237), .B1(n6265), .B2(
        SRAM_192X32_data_out[10]), .O(n2714) );
  INV1S U7173 ( .I(SRAM_192X32_out_decode[1]), .O(n6238) );
  MOAI1S U7174 ( .A1(conv_sram_stop_flag_reg), .A2(n6238), .B1(n6265), .B2(
        SRAM_192X32_data_out[1]), .O(n2713) );
  INV1S U7175 ( .I(SRAM_192X32_out_decode[0]), .O(n6239) );
  MOAI1S U7176 ( .A1(conv_sram_stop_flag_reg), .A2(n6239), .B1(n6265), .B2(
        SRAM_192X32_data_out[0]), .O(n2712) );
  AOI22S U7177 ( .A1(n6243), .A2(n6242), .B1(n6241), .B2(n6240), .O(n6246) );
  OAI22S U7178 ( .A1(n6246), .A2(n6245), .B1(n6244), .B2(n6245), .O(n6266) );
  INV1S U7179 ( .I(SRAM_64X32_out_decode[9]), .O(n6247) );
  MOAI1S U7180 ( .A1(conv_sram_stop_flag_reg), .A2(n6247), .B1(n6265), .B2(
        SRAM_64X32_data_out[9]), .O(n2703) );
  INV1S U7181 ( .I(SRAM_64X32_out_decode[8]), .O(n6248) );
  MOAI1S U7182 ( .A1(conv_sram_stop_flag_reg), .A2(n6248), .B1(n6265), .B2(
        SRAM_64X32_data_out[8]), .O(n2702) );
  INV1S U7183 ( .I(SRAM_64X32_out_decode[5]), .O(n6249) );
  MOAI1S U7184 ( .A1(conv_sram_stop_flag_reg), .A2(n6249), .B1(n6265), .B2(
        SRAM_64X32_data_out[5]), .O(n2699) );
  INV1S U7185 ( .I(SRAM_64X32_out_decode[4]), .O(n6250) );
  MOAI1S U7186 ( .A1(conv_sram_stop_flag_reg), .A2(n6250), .B1(n6265), .B2(
        SRAM_64X32_data_out[4]), .O(n2698) );
  INV1S U7187 ( .I(SRAM_64X32_out_decode[31]), .O(n6251) );
  MOAI1S U7188 ( .A1(conv_sram_stop_flag_reg), .A2(n6251), .B1(n6265), .B2(
        SRAM_64X32_data_out[31]), .O(n2697) );
  INV1S U7189 ( .I(SRAM_64X32_out_decode[30]), .O(n6252) );
  MOAI1S U7190 ( .A1(conv_sram_stop_flag_reg), .A2(n6252), .B1(
        conv_sram_stop_flag_reg), .B2(SRAM_64X32_data_out[30]), .O(n2696) );
  INV1S U7191 ( .I(SRAM_64X32_out_decode[3]), .O(n6253) );
  MOAI1S U7192 ( .A1(conv_sram_stop_flag_reg), .A2(n6253), .B1(n6265), .B2(
        SRAM_64X32_data_out[3]), .O(n2695) );
  INV1S U7193 ( .I(SRAM_64X32_out_decode[29]), .O(n6254) );
  MOAI1S U7194 ( .A1(conv_sram_stop_flag_reg), .A2(n6254), .B1(n6265), .B2(
        SRAM_64X32_data_out[29]), .O(n2694) );
  INV1S U7195 ( .I(SRAM_64X32_out_decode[28]), .O(n6255) );
  MOAI1S U7196 ( .A1(conv_sram_stop_flag_reg), .A2(n6255), .B1(
        conv_sram_stop_flag_reg), .B2(SRAM_64X32_data_out[28]), .O(n2693) );
  INV1S U7197 ( .I(SRAM_64X32_out_decode[27]), .O(n6256) );
  MOAI1S U7198 ( .A1(conv_sram_stop_flag_reg), .A2(n6256), .B1(n6265), .B2(
        SRAM_64X32_data_out[27]), .O(n2692) );
  INV1S U7199 ( .I(SRAM_64X32_out_decode[26]), .O(n6257) );
  MOAI1S U7200 ( .A1(conv_sram_stop_flag_reg), .A2(n6257), .B1(n6265), .B2(
        SRAM_64X32_data_out[26]), .O(n2691) );
  INV1S U7201 ( .I(SRAM_64X32_out_decode[25]), .O(n6258) );
  MOAI1S U7202 ( .A1(conv_sram_stop_flag_reg), .A2(n6258), .B1(n6265), .B2(
        SRAM_64X32_data_out[25]), .O(n2690) );
  INV1S U7203 ( .I(SRAM_64X32_out_decode[24]), .O(n6259) );
  MOAI1S U7204 ( .A1(conv_sram_stop_flag_reg), .A2(n6259), .B1(n6265), .B2(
        SRAM_64X32_data_out[24]), .O(n2689) );
  INV1S U7205 ( .I(SRAM_64X32_out_decode[23]), .O(n6260) );
  MOAI1S U7206 ( .A1(conv_sram_stop_flag_reg), .A2(n6260), .B1(n6265), .B2(
        SRAM_64X32_data_out[23]), .O(n2688) );
  INV1S U7207 ( .I(SRAM_64X32_out_decode[22]), .O(n6261) );
  MOAI1S U7208 ( .A1(conv_sram_stop_flag_reg), .A2(n6261), .B1(n6265), .B2(
        SRAM_64X32_data_out[22]), .O(n2687) );
  INV1S U7209 ( .I(SRAM_64X32_out_decode[21]), .O(n6262) );
  MOAI1S U7210 ( .A1(conv_sram_stop_flag_reg), .A2(n6262), .B1(n6265), .B2(
        SRAM_64X32_data_out[21]), .O(n2686) );
  INV1S U7211 ( .I(SRAM_64X32_out_decode[0]), .O(n6264) );
  MOAI1S U7212 ( .A1(n6265), .A2(n6264), .B1(conv_sram_stop_flag_reg), .B2(
        SRAM_64X32_data_out[0]), .O(n2624) );
  FA1 U7213 ( .A(image[7]), .B(n6271), .CI(n6270), .CO(n6267), .S(n6272) );
  MOAI1S U7214 ( .A1(n3493), .A2(n6273), .B1(n3493), .B2(n6272), .O(n2613) );
  FA1 U7215 ( .A(image[6]), .B(n6275), .CI(n6274), .CO(n6270), .S(n6276) );
  MOAI1S U7216 ( .A1(n3493), .A2(n6277), .B1(n3493), .B2(n6276), .O(n2612) );
  FA1 U7217 ( .A(image[5]), .B(n6279), .CI(n6278), .CO(n6274), .S(n6280) );
  MOAI1S U7218 ( .A1(n3493), .A2(n6281), .B1(n3493), .B2(n6280), .O(n2611) );
  FA1 U7219 ( .A(image[4]), .B(n6283), .CI(n6282), .CO(n6278), .S(n6284) );
  MOAI1S U7220 ( .A1(n3493), .A2(n6285), .B1(n3493), .B2(n6284), .O(n2610) );
  FA1 U7221 ( .A(image[3]), .B(n6287), .CI(n6286), .CO(n6282), .S(n6288) );
  MOAI1S U7222 ( .A1(n3493), .A2(n6289), .B1(n3493), .B2(n6288), .O(n2609) );
  FA1 U7223 ( .A(image[2]), .B(n62910), .CI(n6290), .CO(n6286), .S(n6292) );
  MOAI1S U7224 ( .A1(n3493), .A2(n6293), .B1(n3493), .B2(n6292), .O(n2608) );
  FA1 U7225 ( .A(image[1]), .B(n6295), .CI(n6294), .CO(n6290), .S(n6296) );
  FACS1S U7226 ( .CI1(mult_x_231_n9), .B(mult_x_231_n39), .A(mult_x_231_n48), 
        .CI0(mult_x_231_n10), .CS(mult_x_231_n11), .CO1(mult_x_231_n7), .CO0(
        mult_x_231_n8), .S(N6124) );
endmodule

