# 
#              Synchronous High Speed Single Port SRAM Compiler 
# 
#                    UMC 0.18um GenericII Logic Process
#    __________________________________________________________________________
# 
# 
#      (C) Copyright 2002-2009 Faraday Technology Corp. All Rights Reserved.
#    
#    This source code is an unpublished work belongs to Faraday Technology
#    Corp.  It is considered a trade secret and is not to be divulged or
#    used by parties who have not received written authorization from
#    Faraday Technology Corp.
#    
#    Faraday's home page can be found at:
#    http://www.faraday-tech.com/
#   
#       Module Name      : SRAM_64X32
#       Words            : 64
#       Bits             : 32
#       Byte-Write       : 1
#       Aspect Ratio     : 1
#       Output Loading   : 0.05  (pf)
#       Data Slew        : 0.02  (ns)
#       CK Slew          : 0.02  (ns)
#       Power Ring Width : 2  (um)
# 
# -----------------------------------------------------------------------------
# 
#       Library          : FSA0M_A
#       Memaker          : 200901.2.1
#       Date             : 2024/11/25 18:33:46
# 
# -----------------------------------------------------------------------------


NAMESCASESENSITIVE ON ;
MACRO SRAM_64X32
CLASS BLOCK ;
FOREIGN SRAM_64X32 0.000 0.000 ;
ORIGIN 0.000 0.000 ;
SIZE 531.960 BY 156.800 ;
SYMMETRY x y r90 ;
SITE core ;
PIN GND
  DIRECTION INOUT ;
  USE GROUND ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 530.840 129.700 531.960 132.940 ;
  LAYER ME3 ;
  RECT 530.840 129.700 531.960 132.940 ;
  LAYER ME2 ;
  RECT 530.840 129.700 531.960 132.940 ;
  LAYER ME1 ;
  RECT 530.840 129.700 531.960 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 121.860 531.960 125.100 ;
  LAYER ME3 ;
  RECT 530.840 121.860 531.960 125.100 ;
  LAYER ME2 ;
  RECT 530.840 121.860 531.960 125.100 ;
  LAYER ME1 ;
  RECT 530.840 121.860 531.960 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 114.020 531.960 117.260 ;
  LAYER ME3 ;
  RECT 530.840 114.020 531.960 117.260 ;
  LAYER ME2 ;
  RECT 530.840 114.020 531.960 117.260 ;
  LAYER ME1 ;
  RECT 530.840 114.020 531.960 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 106.180 531.960 109.420 ;
  LAYER ME3 ;
  RECT 530.840 106.180 531.960 109.420 ;
  LAYER ME2 ;
  RECT 530.840 106.180 531.960 109.420 ;
  LAYER ME1 ;
  RECT 530.840 106.180 531.960 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 98.340 531.960 101.580 ;
  LAYER ME3 ;
  RECT 530.840 98.340 531.960 101.580 ;
  LAYER ME2 ;
  RECT 530.840 98.340 531.960 101.580 ;
  LAYER ME1 ;
  RECT 530.840 98.340 531.960 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 90.500 531.960 93.740 ;
  LAYER ME3 ;
  RECT 530.840 90.500 531.960 93.740 ;
  LAYER ME2 ;
  RECT 530.840 90.500 531.960 93.740 ;
  LAYER ME1 ;
  RECT 530.840 90.500 531.960 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 51.300 531.960 54.540 ;
  LAYER ME3 ;
  RECT 530.840 51.300 531.960 54.540 ;
  LAYER ME2 ;
  RECT 530.840 51.300 531.960 54.540 ;
  LAYER ME1 ;
  RECT 530.840 51.300 531.960 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 43.460 531.960 46.700 ;
  LAYER ME3 ;
  RECT 530.840 43.460 531.960 46.700 ;
  LAYER ME2 ;
  RECT 530.840 43.460 531.960 46.700 ;
  LAYER ME1 ;
  RECT 530.840 43.460 531.960 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 35.620 531.960 38.860 ;
  LAYER ME3 ;
  RECT 530.840 35.620 531.960 38.860 ;
  LAYER ME2 ;
  RECT 530.840 35.620 531.960 38.860 ;
  LAYER ME1 ;
  RECT 530.840 35.620 531.960 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 27.780 531.960 31.020 ;
  LAYER ME3 ;
  RECT 530.840 27.780 531.960 31.020 ;
  LAYER ME2 ;
  RECT 530.840 27.780 531.960 31.020 ;
  LAYER ME1 ;
  RECT 530.840 27.780 531.960 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 19.940 531.960 23.180 ;
  LAYER ME3 ;
  RECT 530.840 19.940 531.960 23.180 ;
  LAYER ME2 ;
  RECT 530.840 19.940 531.960 23.180 ;
  LAYER ME1 ;
  RECT 530.840 19.940 531.960 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 12.100 531.960 15.340 ;
  LAYER ME3 ;
  RECT 530.840 12.100 531.960 15.340 ;
  LAYER ME2 ;
  RECT 530.840 12.100 531.960 15.340 ;
  LAYER ME1 ;
  RECT 530.840 12.100 531.960 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME3 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME2 ;
  RECT 0.000 129.700 1.120 132.940 ;
  LAYER ME1 ;
  RECT 0.000 129.700 1.120 132.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME3 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME2 ;
  RECT 0.000 121.860 1.120 125.100 ;
  LAYER ME1 ;
  RECT 0.000 121.860 1.120 125.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME3 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME2 ;
  RECT 0.000 114.020 1.120 117.260 ;
  LAYER ME1 ;
  RECT 0.000 114.020 1.120 117.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME3 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME2 ;
  RECT 0.000 106.180 1.120 109.420 ;
  LAYER ME1 ;
  RECT 0.000 106.180 1.120 109.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME3 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME2 ;
  RECT 0.000 98.340 1.120 101.580 ;
  LAYER ME1 ;
  RECT 0.000 98.340 1.120 101.580 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME3 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME2 ;
  RECT 0.000 90.500 1.120 93.740 ;
  LAYER ME1 ;
  RECT 0.000 90.500 1.120 93.740 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME3 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME2 ;
  RECT 0.000 51.300 1.120 54.540 ;
  LAYER ME1 ;
  RECT 0.000 51.300 1.120 54.540 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME3 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME2 ;
  RECT 0.000 43.460 1.120 46.700 ;
  LAYER ME1 ;
  RECT 0.000 43.460 1.120 46.700 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME3 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME2 ;
  RECT 0.000 35.620 1.120 38.860 ;
  LAYER ME1 ;
  RECT 0.000 35.620 1.120 38.860 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME3 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME2 ;
  RECT 0.000 27.780 1.120 31.020 ;
  LAYER ME1 ;
  RECT 0.000 27.780 1.120 31.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME3 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME2 ;
  RECT 0.000 19.940 1.120 23.180 ;
  LAYER ME1 ;
  RECT 0.000 19.940 1.120 23.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME3 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME2 ;
  RECT 0.000 12.100 1.120 15.340 ;
  LAYER ME1 ;
  RECT 0.000 12.100 1.120 15.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 489.580 155.680 493.120 156.800 ;
  LAYER ME3 ;
  RECT 489.580 155.680 493.120 156.800 ;
  LAYER ME2 ;
  RECT 489.580 155.680 493.120 156.800 ;
  LAYER ME1 ;
  RECT 489.580 155.680 493.120 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 480.900 155.680 484.440 156.800 ;
  LAYER ME3 ;
  RECT 480.900 155.680 484.440 156.800 ;
  LAYER ME2 ;
  RECT 480.900 155.680 484.440 156.800 ;
  LAYER ME1 ;
  RECT 480.900 155.680 484.440 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 472.220 155.680 475.760 156.800 ;
  LAYER ME3 ;
  RECT 472.220 155.680 475.760 156.800 ;
  LAYER ME2 ;
  RECT 472.220 155.680 475.760 156.800 ;
  LAYER ME1 ;
  RECT 472.220 155.680 475.760 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 463.540 155.680 467.080 156.800 ;
  LAYER ME3 ;
  RECT 463.540 155.680 467.080 156.800 ;
  LAYER ME2 ;
  RECT 463.540 155.680 467.080 156.800 ;
  LAYER ME1 ;
  RECT 463.540 155.680 467.080 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 454.860 155.680 458.400 156.800 ;
  LAYER ME3 ;
  RECT 454.860 155.680 458.400 156.800 ;
  LAYER ME2 ;
  RECT 454.860 155.680 458.400 156.800 ;
  LAYER ME1 ;
  RECT 454.860 155.680 458.400 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 446.180 155.680 449.720 156.800 ;
  LAYER ME3 ;
  RECT 446.180 155.680 449.720 156.800 ;
  LAYER ME2 ;
  RECT 446.180 155.680 449.720 156.800 ;
  LAYER ME1 ;
  RECT 446.180 155.680 449.720 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 402.780 155.680 406.320 156.800 ;
  LAYER ME3 ;
  RECT 402.780 155.680 406.320 156.800 ;
  LAYER ME2 ;
  RECT 402.780 155.680 406.320 156.800 ;
  LAYER ME1 ;
  RECT 402.780 155.680 406.320 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 394.100 155.680 397.640 156.800 ;
  LAYER ME3 ;
  RECT 394.100 155.680 397.640 156.800 ;
  LAYER ME2 ;
  RECT 394.100 155.680 397.640 156.800 ;
  LAYER ME1 ;
  RECT 394.100 155.680 397.640 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 385.420 155.680 388.960 156.800 ;
  LAYER ME3 ;
  RECT 385.420 155.680 388.960 156.800 ;
  LAYER ME2 ;
  RECT 385.420 155.680 388.960 156.800 ;
  LAYER ME1 ;
  RECT 385.420 155.680 388.960 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 376.740 155.680 380.280 156.800 ;
  LAYER ME3 ;
  RECT 376.740 155.680 380.280 156.800 ;
  LAYER ME2 ;
  RECT 376.740 155.680 380.280 156.800 ;
  LAYER ME1 ;
  RECT 376.740 155.680 380.280 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 368.060 155.680 371.600 156.800 ;
  LAYER ME3 ;
  RECT 368.060 155.680 371.600 156.800 ;
  LAYER ME2 ;
  RECT 368.060 155.680 371.600 156.800 ;
  LAYER ME1 ;
  RECT 368.060 155.680 371.600 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 359.380 155.680 362.920 156.800 ;
  LAYER ME3 ;
  RECT 359.380 155.680 362.920 156.800 ;
  LAYER ME2 ;
  RECT 359.380 155.680 362.920 156.800 ;
  LAYER ME1 ;
  RECT 359.380 155.680 362.920 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 315.980 155.680 319.520 156.800 ;
  LAYER ME3 ;
  RECT 315.980 155.680 319.520 156.800 ;
  LAYER ME2 ;
  RECT 315.980 155.680 319.520 156.800 ;
  LAYER ME1 ;
  RECT 315.980 155.680 319.520 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 307.300 155.680 310.840 156.800 ;
  LAYER ME3 ;
  RECT 307.300 155.680 310.840 156.800 ;
  LAYER ME2 ;
  RECT 307.300 155.680 310.840 156.800 ;
  LAYER ME1 ;
  RECT 307.300 155.680 310.840 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 298.620 155.680 302.160 156.800 ;
  LAYER ME3 ;
  RECT 298.620 155.680 302.160 156.800 ;
  LAYER ME2 ;
  RECT 298.620 155.680 302.160 156.800 ;
  LAYER ME1 ;
  RECT 298.620 155.680 302.160 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER ME3 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER ME2 ;
  RECT 289.940 155.680 293.480 156.800 ;
  LAYER ME1 ;
  RECT 289.940 155.680 293.480 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER ME3 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER ME2 ;
  RECT 281.260 155.680 284.800 156.800 ;
  LAYER ME1 ;
  RECT 281.260 155.680 284.800 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER ME3 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER ME2 ;
  RECT 272.580 155.680 276.120 156.800 ;
  LAYER ME1 ;
  RECT 272.580 155.680 276.120 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER ME3 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER ME2 ;
  RECT 229.180 155.680 232.720 156.800 ;
  LAYER ME1 ;
  RECT 229.180 155.680 232.720 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER ME3 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER ME2 ;
  RECT 220.500 155.680 224.040 156.800 ;
  LAYER ME1 ;
  RECT 220.500 155.680 224.040 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER ME3 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER ME2 ;
  RECT 211.820 155.680 215.360 156.800 ;
  LAYER ME1 ;
  RECT 211.820 155.680 215.360 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER ME3 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER ME2 ;
  RECT 203.140 155.680 206.680 156.800 ;
  LAYER ME1 ;
  RECT 203.140 155.680 206.680 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER ME3 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER ME2 ;
  RECT 194.460 155.680 198.000 156.800 ;
  LAYER ME1 ;
  RECT 194.460 155.680 198.000 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER ME3 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER ME2 ;
  RECT 185.780 155.680 189.320 156.800 ;
  LAYER ME1 ;
  RECT 185.780 155.680 189.320 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER ME3 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER ME2 ;
  RECT 142.380 155.680 145.920 156.800 ;
  LAYER ME1 ;
  RECT 142.380 155.680 145.920 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER ME3 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER ME2 ;
  RECT 133.700 155.680 137.240 156.800 ;
  LAYER ME1 ;
  RECT 133.700 155.680 137.240 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER ME3 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER ME2 ;
  RECT 125.020 155.680 128.560 156.800 ;
  LAYER ME1 ;
  RECT 125.020 155.680 128.560 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER ME3 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER ME2 ;
  RECT 116.340 155.680 119.880 156.800 ;
  LAYER ME1 ;
  RECT 116.340 155.680 119.880 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER ME3 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER ME2 ;
  RECT 107.660 155.680 111.200 156.800 ;
  LAYER ME1 ;
  RECT 107.660 155.680 111.200 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER ME3 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER ME2 ;
  RECT 98.980 155.680 102.520 156.800 ;
  LAYER ME1 ;
  RECT 98.980 155.680 102.520 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER ME3 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER ME2 ;
  RECT 55.580 155.680 59.120 156.800 ;
  LAYER ME1 ;
  RECT 55.580 155.680 59.120 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER ME3 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER ME2 ;
  RECT 46.900 155.680 50.440 156.800 ;
  LAYER ME1 ;
  RECT 46.900 155.680 50.440 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER ME3 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER ME2 ;
  RECT 38.220 155.680 41.760 156.800 ;
  LAYER ME1 ;
  RECT 38.220 155.680 41.760 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER ME3 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER ME2 ;
  RECT 29.540 155.680 33.080 156.800 ;
  LAYER ME1 ;
  RECT 29.540 155.680 33.080 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER ME3 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER ME2 ;
  RECT 20.860 155.680 24.400 156.800 ;
  LAYER ME1 ;
  RECT 20.860 155.680 24.400 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER ME3 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER ME2 ;
  RECT 12.180 155.680 15.720 156.800 ;
  LAYER ME1 ;
  RECT 12.180 155.680 15.720 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER ME3 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER ME2 ;
  RECT 511.900 0.000 515.440 1.120 ;
  LAYER ME1 ;
  RECT 511.900 0.000 515.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER ME3 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER ME2 ;
  RECT 490.200 0.000 493.740 1.120 ;
  LAYER ME1 ;
  RECT 490.200 0.000 493.740 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME3 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME2 ;
  RECT 468.500 0.000 472.040 1.120 ;
  LAYER ME1 ;
  RECT 468.500 0.000 472.040 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.660 0.000 359.200 1.120 ;
  LAYER ME3 ;
  RECT 355.660 0.000 359.200 1.120 ;
  LAYER ME2 ;
  RECT 355.660 0.000 359.200 1.120 ;
  LAYER ME1 ;
  RECT 355.660 0.000 359.200 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 329.000 0.000 332.540 1.120 ;
  LAYER ME3 ;
  RECT 329.000 0.000 332.540 1.120 ;
  LAYER ME2 ;
  RECT 329.000 0.000 332.540 1.120 ;
  LAYER ME1 ;
  RECT 329.000 0.000 332.540 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 312.260 0.000 315.800 1.120 ;
  LAYER ME3 ;
  RECT 312.260 0.000 315.800 1.120 ;
  LAYER ME2 ;
  RECT 312.260 0.000 315.800 1.120 ;
  LAYER ME1 ;
  RECT 312.260 0.000 315.800 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.300 0.000 279.840 1.120 ;
  LAYER ME3 ;
  RECT 276.300 0.000 279.840 1.120 ;
  LAYER ME2 ;
  RECT 276.300 0.000 279.840 1.120 ;
  LAYER ME1 ;
  RECT 276.300 0.000 279.840 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER ME3 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER ME2 ;
  RECT 267.620 0.000 271.160 1.120 ;
  LAYER ME1 ;
  RECT 267.620 0.000 271.160 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME3 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME2 ;
  RECT 246.540 0.000 250.080 1.120 ;
  LAYER ME1 ;
  RECT 246.540 0.000 250.080 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME3 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME2 ;
  RECT 139.900 0.000 143.440 1.120 ;
  LAYER ME1 ;
  RECT 139.900 0.000 143.440 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME3 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME2 ;
  RECT 113.860 0.000 117.400 1.120 ;
  LAYER ME1 ;
  RECT 113.860 0.000 117.400 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME3 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME2 ;
  RECT 92.160 0.000 95.700 1.120 ;
  LAYER ME1 ;
  RECT 92.160 0.000 95.700 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME3 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME2 ;
  RECT 70.460 0.000 74.000 1.120 ;
  LAYER ME1 ;
  RECT 70.460 0.000 74.000 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME3 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME2 ;
  RECT 43.800 0.000 47.340 1.120 ;
  LAYER ME1 ;
  RECT 43.800 0.000 47.340 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME3 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME2 ;
  RECT 27.060 0.000 30.600 1.120 ;
  LAYER ME1 ;
  RECT 27.060 0.000 30.600 1.120 ;
 END
END GND
PIN VCC
  DIRECTION INOUT ;
  USE POWER ;
  SHAPE ABUTMENT ;
 PORT
  LAYER ME4 ;
  RECT 530.840 125.780 531.960 129.020 ;
  LAYER ME3 ;
  RECT 530.840 125.780 531.960 129.020 ;
  LAYER ME2 ;
  RECT 530.840 125.780 531.960 129.020 ;
  LAYER ME1 ;
  RECT 530.840 125.780 531.960 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 117.940 531.960 121.180 ;
  LAYER ME3 ;
  RECT 530.840 117.940 531.960 121.180 ;
  LAYER ME2 ;
  RECT 530.840 117.940 531.960 121.180 ;
  LAYER ME1 ;
  RECT 530.840 117.940 531.960 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 110.100 531.960 113.340 ;
  LAYER ME3 ;
  RECT 530.840 110.100 531.960 113.340 ;
  LAYER ME2 ;
  RECT 530.840 110.100 531.960 113.340 ;
  LAYER ME1 ;
  RECT 530.840 110.100 531.960 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 102.260 531.960 105.500 ;
  LAYER ME3 ;
  RECT 530.840 102.260 531.960 105.500 ;
  LAYER ME2 ;
  RECT 530.840 102.260 531.960 105.500 ;
  LAYER ME1 ;
  RECT 530.840 102.260 531.960 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 94.420 531.960 97.660 ;
  LAYER ME3 ;
  RECT 530.840 94.420 531.960 97.660 ;
  LAYER ME2 ;
  RECT 530.840 94.420 531.960 97.660 ;
  LAYER ME1 ;
  RECT 530.840 94.420 531.960 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 86.580 531.960 89.820 ;
  LAYER ME3 ;
  RECT 530.840 86.580 531.960 89.820 ;
  LAYER ME2 ;
  RECT 530.840 86.580 531.960 89.820 ;
  LAYER ME1 ;
  RECT 530.840 86.580 531.960 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 47.380 531.960 50.620 ;
  LAYER ME3 ;
  RECT 530.840 47.380 531.960 50.620 ;
  LAYER ME2 ;
  RECT 530.840 47.380 531.960 50.620 ;
  LAYER ME1 ;
  RECT 530.840 47.380 531.960 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 39.540 531.960 42.780 ;
  LAYER ME3 ;
  RECT 530.840 39.540 531.960 42.780 ;
  LAYER ME2 ;
  RECT 530.840 39.540 531.960 42.780 ;
  LAYER ME1 ;
  RECT 530.840 39.540 531.960 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 31.700 531.960 34.940 ;
  LAYER ME3 ;
  RECT 530.840 31.700 531.960 34.940 ;
  LAYER ME2 ;
  RECT 530.840 31.700 531.960 34.940 ;
  LAYER ME1 ;
  RECT 530.840 31.700 531.960 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 23.860 531.960 27.100 ;
  LAYER ME3 ;
  RECT 530.840 23.860 531.960 27.100 ;
  LAYER ME2 ;
  RECT 530.840 23.860 531.960 27.100 ;
  LAYER ME1 ;
  RECT 530.840 23.860 531.960 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 16.020 531.960 19.260 ;
  LAYER ME3 ;
  RECT 530.840 16.020 531.960 19.260 ;
  LAYER ME2 ;
  RECT 530.840 16.020 531.960 19.260 ;
  LAYER ME1 ;
  RECT 530.840 16.020 531.960 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 530.840 8.180 531.960 11.420 ;
  LAYER ME3 ;
  RECT 530.840 8.180 531.960 11.420 ;
  LAYER ME2 ;
  RECT 530.840 8.180 531.960 11.420 ;
  LAYER ME1 ;
  RECT 530.840 8.180 531.960 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME3 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME2 ;
  RECT 0.000 125.780 1.120 129.020 ;
  LAYER ME1 ;
  RECT 0.000 125.780 1.120 129.020 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME3 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME2 ;
  RECT 0.000 117.940 1.120 121.180 ;
  LAYER ME1 ;
  RECT 0.000 117.940 1.120 121.180 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME3 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME2 ;
  RECT 0.000 110.100 1.120 113.340 ;
  LAYER ME1 ;
  RECT 0.000 110.100 1.120 113.340 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME3 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME2 ;
  RECT 0.000 102.260 1.120 105.500 ;
  LAYER ME1 ;
  RECT 0.000 102.260 1.120 105.500 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME3 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME2 ;
  RECT 0.000 94.420 1.120 97.660 ;
  LAYER ME1 ;
  RECT 0.000 94.420 1.120 97.660 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME3 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME2 ;
  RECT 0.000 86.580 1.120 89.820 ;
  LAYER ME1 ;
  RECT 0.000 86.580 1.120 89.820 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME3 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME2 ;
  RECT 0.000 47.380 1.120 50.620 ;
  LAYER ME1 ;
  RECT 0.000 47.380 1.120 50.620 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME3 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME2 ;
  RECT 0.000 39.540 1.120 42.780 ;
  LAYER ME1 ;
  RECT 0.000 39.540 1.120 42.780 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME3 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME2 ;
  RECT 0.000 31.700 1.120 34.940 ;
  LAYER ME1 ;
  RECT 0.000 31.700 1.120 34.940 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME3 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME2 ;
  RECT 0.000 23.860 1.120 27.100 ;
  LAYER ME1 ;
  RECT 0.000 23.860 1.120 27.100 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME3 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME2 ;
  RECT 0.000 16.020 1.120 19.260 ;
  LAYER ME1 ;
  RECT 0.000 16.020 1.120 19.260 ;
 END
 PORT
  LAYER ME4 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME3 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME2 ;
  RECT 0.000 8.180 1.120 11.420 ;
  LAYER ME1 ;
  RECT 0.000 8.180 1.120 11.420 ;
 END
 PORT
  LAYER ME4 ;
  RECT 485.240 155.680 488.780 156.800 ;
  LAYER ME3 ;
  RECT 485.240 155.680 488.780 156.800 ;
  LAYER ME2 ;
  RECT 485.240 155.680 488.780 156.800 ;
  LAYER ME1 ;
  RECT 485.240 155.680 488.780 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 476.560 155.680 480.100 156.800 ;
  LAYER ME3 ;
  RECT 476.560 155.680 480.100 156.800 ;
  LAYER ME2 ;
  RECT 476.560 155.680 480.100 156.800 ;
  LAYER ME1 ;
  RECT 476.560 155.680 480.100 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 467.880 155.680 471.420 156.800 ;
  LAYER ME3 ;
  RECT 467.880 155.680 471.420 156.800 ;
  LAYER ME2 ;
  RECT 467.880 155.680 471.420 156.800 ;
  LAYER ME1 ;
  RECT 467.880 155.680 471.420 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 459.200 155.680 462.740 156.800 ;
  LAYER ME3 ;
  RECT 459.200 155.680 462.740 156.800 ;
  LAYER ME2 ;
  RECT 459.200 155.680 462.740 156.800 ;
  LAYER ME1 ;
  RECT 459.200 155.680 462.740 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 450.520 155.680 454.060 156.800 ;
  LAYER ME3 ;
  RECT 450.520 155.680 454.060 156.800 ;
  LAYER ME2 ;
  RECT 450.520 155.680 454.060 156.800 ;
  LAYER ME1 ;
  RECT 450.520 155.680 454.060 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 441.840 155.680 445.380 156.800 ;
  LAYER ME3 ;
  RECT 441.840 155.680 445.380 156.800 ;
  LAYER ME2 ;
  RECT 441.840 155.680 445.380 156.800 ;
  LAYER ME1 ;
  RECT 441.840 155.680 445.380 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 398.440 155.680 401.980 156.800 ;
  LAYER ME3 ;
  RECT 398.440 155.680 401.980 156.800 ;
  LAYER ME2 ;
  RECT 398.440 155.680 401.980 156.800 ;
  LAYER ME1 ;
  RECT 398.440 155.680 401.980 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 389.760 155.680 393.300 156.800 ;
  LAYER ME3 ;
  RECT 389.760 155.680 393.300 156.800 ;
  LAYER ME2 ;
  RECT 389.760 155.680 393.300 156.800 ;
  LAYER ME1 ;
  RECT 389.760 155.680 393.300 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 381.080 155.680 384.620 156.800 ;
  LAYER ME3 ;
  RECT 381.080 155.680 384.620 156.800 ;
  LAYER ME2 ;
  RECT 381.080 155.680 384.620 156.800 ;
  LAYER ME1 ;
  RECT 381.080 155.680 384.620 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 372.400 155.680 375.940 156.800 ;
  LAYER ME3 ;
  RECT 372.400 155.680 375.940 156.800 ;
  LAYER ME2 ;
  RECT 372.400 155.680 375.940 156.800 ;
  LAYER ME1 ;
  RECT 372.400 155.680 375.940 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 363.720 155.680 367.260 156.800 ;
  LAYER ME3 ;
  RECT 363.720 155.680 367.260 156.800 ;
  LAYER ME2 ;
  RECT 363.720 155.680 367.260 156.800 ;
  LAYER ME1 ;
  RECT 363.720 155.680 367.260 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 355.040 155.680 358.580 156.800 ;
  LAYER ME3 ;
  RECT 355.040 155.680 358.580 156.800 ;
  LAYER ME2 ;
  RECT 355.040 155.680 358.580 156.800 ;
  LAYER ME1 ;
  RECT 355.040 155.680 358.580 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 311.640 155.680 315.180 156.800 ;
  LAYER ME3 ;
  RECT 311.640 155.680 315.180 156.800 ;
  LAYER ME2 ;
  RECT 311.640 155.680 315.180 156.800 ;
  LAYER ME1 ;
  RECT 311.640 155.680 315.180 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 302.960 155.680 306.500 156.800 ;
  LAYER ME3 ;
  RECT 302.960 155.680 306.500 156.800 ;
  LAYER ME2 ;
  RECT 302.960 155.680 306.500 156.800 ;
  LAYER ME1 ;
  RECT 302.960 155.680 306.500 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER ME3 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER ME2 ;
  RECT 294.280 155.680 297.820 156.800 ;
  LAYER ME1 ;
  RECT 294.280 155.680 297.820 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER ME3 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER ME2 ;
  RECT 285.600 155.680 289.140 156.800 ;
  LAYER ME1 ;
  RECT 285.600 155.680 289.140 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER ME3 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER ME2 ;
  RECT 276.920 155.680 280.460 156.800 ;
  LAYER ME1 ;
  RECT 276.920 155.680 280.460 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER ME3 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER ME2 ;
  RECT 268.240 155.680 271.780 156.800 ;
  LAYER ME1 ;
  RECT 268.240 155.680 271.780 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER ME3 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER ME2 ;
  RECT 224.840 155.680 228.380 156.800 ;
  LAYER ME1 ;
  RECT 224.840 155.680 228.380 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER ME3 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER ME2 ;
  RECT 216.160 155.680 219.700 156.800 ;
  LAYER ME1 ;
  RECT 216.160 155.680 219.700 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER ME3 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER ME2 ;
  RECT 207.480 155.680 211.020 156.800 ;
  LAYER ME1 ;
  RECT 207.480 155.680 211.020 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER ME3 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER ME2 ;
  RECT 198.800 155.680 202.340 156.800 ;
  LAYER ME1 ;
  RECT 198.800 155.680 202.340 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER ME3 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER ME2 ;
  RECT 190.120 155.680 193.660 156.800 ;
  LAYER ME1 ;
  RECT 190.120 155.680 193.660 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER ME3 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER ME2 ;
  RECT 181.440 155.680 184.980 156.800 ;
  LAYER ME1 ;
  RECT 181.440 155.680 184.980 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER ME3 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER ME2 ;
  RECT 138.040 155.680 141.580 156.800 ;
  LAYER ME1 ;
  RECT 138.040 155.680 141.580 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER ME3 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER ME2 ;
  RECT 129.360 155.680 132.900 156.800 ;
  LAYER ME1 ;
  RECT 129.360 155.680 132.900 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER ME3 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER ME2 ;
  RECT 120.680 155.680 124.220 156.800 ;
  LAYER ME1 ;
  RECT 120.680 155.680 124.220 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER ME3 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER ME2 ;
  RECT 112.000 155.680 115.540 156.800 ;
  LAYER ME1 ;
  RECT 112.000 155.680 115.540 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER ME3 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER ME2 ;
  RECT 103.320 155.680 106.860 156.800 ;
  LAYER ME1 ;
  RECT 103.320 155.680 106.860 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER ME3 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER ME2 ;
  RECT 94.640 155.680 98.180 156.800 ;
  LAYER ME1 ;
  RECT 94.640 155.680 98.180 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER ME3 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER ME2 ;
  RECT 51.240 155.680 54.780 156.800 ;
  LAYER ME1 ;
  RECT 51.240 155.680 54.780 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER ME3 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER ME2 ;
  RECT 42.560 155.680 46.100 156.800 ;
  LAYER ME1 ;
  RECT 42.560 155.680 46.100 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER ME3 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER ME2 ;
  RECT 33.880 155.680 37.420 156.800 ;
  LAYER ME1 ;
  RECT 33.880 155.680 37.420 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER ME3 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER ME2 ;
  RECT 25.200 155.680 28.740 156.800 ;
  LAYER ME1 ;
  RECT 25.200 155.680 28.740 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER ME3 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER ME2 ;
  RECT 16.520 155.680 20.060 156.800 ;
  LAYER ME1 ;
  RECT 16.520 155.680 20.060 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER ME3 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER ME2 ;
  RECT 7.840 155.680 11.380 156.800 ;
  LAYER ME1 ;
  RECT 7.840 155.680 11.380 156.800 ;
 END
 PORT
  LAYER ME4 ;
  RECT 520.580 0.000 524.120 1.120 ;
  LAYER ME3 ;
  RECT 520.580 0.000 524.120 1.120 ;
  LAYER ME2 ;
  RECT 520.580 0.000 524.120 1.120 ;
  LAYER ME1 ;
  RECT 520.580 0.000 524.120 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 498.880 0.000 502.420 1.120 ;
  LAYER ME3 ;
  RECT 498.880 0.000 502.420 1.120 ;
  LAYER ME2 ;
  RECT 498.880 0.000 502.420 1.120 ;
  LAYER ME1 ;
  RECT 498.880 0.000 502.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 482.140 0.000 485.680 1.120 ;
  LAYER ME3 ;
  RECT 482.140 0.000 485.680 1.120 ;
  LAYER ME2 ;
  RECT 482.140 0.000 485.680 1.120 ;
  LAYER ME1 ;
  RECT 482.140 0.000 485.680 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 455.480 0.000 459.020 1.120 ;
  LAYER ME3 ;
  RECT 455.480 0.000 459.020 1.120 ;
  LAYER ME2 ;
  RECT 455.480 0.000 459.020 1.120 ;
  LAYER ME1 ;
  RECT 455.480 0.000 459.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 342.640 0.000 346.180 1.120 ;
  LAYER ME3 ;
  RECT 342.640 0.000 346.180 1.120 ;
  LAYER ME2 ;
  RECT 342.640 0.000 346.180 1.120 ;
  LAYER ME1 ;
  RECT 342.640 0.000 346.180 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 320.940 0.000 324.480 1.120 ;
  LAYER ME3 ;
  RECT 320.940 0.000 324.480 1.120 ;
  LAYER ME2 ;
  RECT 320.940 0.000 324.480 1.120 ;
  LAYER ME1 ;
  RECT 320.940 0.000 324.480 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 299.240 0.000 302.780 1.120 ;
  LAYER ME3 ;
  RECT 299.240 0.000 302.780 1.120 ;
  LAYER ME2 ;
  RECT 299.240 0.000 302.780 1.120 ;
  LAYER ME1 ;
  RECT 299.240 0.000 302.780 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 271.960 0.000 275.500 1.120 ;
  LAYER ME3 ;
  RECT 271.960 0.000 275.500 1.120 ;
  LAYER ME2 ;
  RECT 271.960 0.000 275.500 1.120 ;
  LAYER ME1 ;
  RECT 271.960 0.000 275.500 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 263.280 0.000 266.820 1.120 ;
  LAYER ME3 ;
  RECT 263.280 0.000 266.820 1.120 ;
  LAYER ME2 ;
  RECT 263.280 0.000 266.820 1.120 ;
  LAYER ME1 ;
  RECT 263.280 0.000 266.820 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER ME3 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER ME2 ;
  RECT 235.380 0.000 238.920 1.120 ;
  LAYER ME1 ;
  RECT 235.380 0.000 238.920 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME3 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME2 ;
  RECT 126.880 0.000 130.420 1.120 ;
  LAYER ME1 ;
  RECT 126.880 0.000 130.420 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME3 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME2 ;
  RECT 100.220 0.000 103.760 1.120 ;
  LAYER ME1 ;
  RECT 100.220 0.000 103.760 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME3 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME2 ;
  RECT 83.480 0.000 87.020 1.120 ;
  LAYER ME1 ;
  RECT 83.480 0.000 87.020 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME3 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME2 ;
  RECT 56.820 0.000 60.360 1.120 ;
  LAYER ME1 ;
  RECT 56.820 0.000 60.360 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME3 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME2 ;
  RECT 35.740 0.000 39.280 1.120 ;
  LAYER ME1 ;
  RECT 35.740 0.000 39.280 1.120 ;
 END
 PORT
  LAYER ME4 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME3 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME2 ;
  RECT 14.040 0.000 17.580 1.120 ;
  LAYER ME1 ;
  RECT 14.040 0.000 17.580 1.120 ;
 END
END VCC
PIN DO31
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 518.380 0.000 519.500 1.120 ;
  LAYER ME3 ;
  RECT 518.380 0.000 519.500 1.120 ;
  LAYER ME2 ;
  RECT 518.380 0.000 519.500 1.120 ;
  LAYER ME1 ;
  RECT 518.380 0.000 519.500 1.120 ;
 END
END DO31
PIN DI31
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME3 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME2 ;
  RECT 509.700 0.000 510.820 1.120 ;
  LAYER ME1 ;
  RECT 509.700 0.000 510.820 1.120 ;
 END
END DI31
PIN DO30
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER ME3 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER ME2 ;
  RECT 504.740 0.000 505.860 1.120 ;
  LAYER ME1 ;
  RECT 504.740 0.000 505.860 1.120 ;
 END
END DO30
PIN DI30
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER ME3 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER ME2 ;
  RECT 496.680 0.000 497.800 1.120 ;
  LAYER ME1 ;
  RECT 496.680 0.000 497.800 1.120 ;
 END
END DI30
PIN DO29
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME3 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME2 ;
  RECT 488.000 0.000 489.120 1.120 ;
  LAYER ME1 ;
  RECT 488.000 0.000 489.120 1.120 ;
 END
END DO29
PIN DI29
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER ME3 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER ME2 ;
  RECT 479.940 0.000 481.060 1.120 ;
  LAYER ME1 ;
  RECT 479.940 0.000 481.060 1.120 ;
 END
END DI29
PIN DO28
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 474.980 0.000 476.100 1.120 ;
  LAYER ME3 ;
  RECT 474.980 0.000 476.100 1.120 ;
  LAYER ME2 ;
  RECT 474.980 0.000 476.100 1.120 ;
  LAYER ME1 ;
  RECT 474.980 0.000 476.100 1.120 ;
 END
END DO28
PIN DI28
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 466.300 0.000 467.420 1.120 ;
  LAYER ME3 ;
  RECT 466.300 0.000 467.420 1.120 ;
  LAYER ME2 ;
  RECT 466.300 0.000 467.420 1.120 ;
  LAYER ME1 ;
  RECT 466.300 0.000 467.420 1.120 ;
 END
END DI28
PIN DO27
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 461.960 0.000 463.080 1.120 ;
  LAYER ME3 ;
  RECT 461.960 0.000 463.080 1.120 ;
  LAYER ME2 ;
  RECT 461.960 0.000 463.080 1.120 ;
  LAYER ME1 ;
  RECT 461.960 0.000 463.080 1.120 ;
 END
END DO27
PIN DI27
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 453.280 0.000 454.400 1.120 ;
  LAYER ME3 ;
  RECT 453.280 0.000 454.400 1.120 ;
  LAYER ME2 ;
  RECT 453.280 0.000 454.400 1.120 ;
  LAYER ME1 ;
  RECT 453.280 0.000 454.400 1.120 ;
 END
END DI27
PIN DO26
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 448.320 0.000 449.440 1.120 ;
  LAYER ME3 ;
  RECT 448.320 0.000 449.440 1.120 ;
  LAYER ME2 ;
  RECT 448.320 0.000 449.440 1.120 ;
  LAYER ME1 ;
  RECT 448.320 0.000 449.440 1.120 ;
 END
END DO26
PIN DI26
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 440.260 0.000 441.380 1.120 ;
  LAYER ME3 ;
  RECT 440.260 0.000 441.380 1.120 ;
  LAYER ME2 ;
  RECT 440.260 0.000 441.380 1.120 ;
  LAYER ME1 ;
  RECT 440.260 0.000 441.380 1.120 ;
 END
END DI26
PIN DO25
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 431.580 0.000 432.700 1.120 ;
  LAYER ME3 ;
  RECT 431.580 0.000 432.700 1.120 ;
  LAYER ME2 ;
  RECT 431.580 0.000 432.700 1.120 ;
  LAYER ME1 ;
  RECT 431.580 0.000 432.700 1.120 ;
 END
END DO25
PIN DI25
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER ME3 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER ME2 ;
  RECT 423.520 0.000 424.640 1.120 ;
  LAYER ME1 ;
  RECT 423.520 0.000 424.640 1.120 ;
 END
END DI25
PIN DO24
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 418.560 0.000 419.680 1.120 ;
  LAYER ME3 ;
  RECT 418.560 0.000 419.680 1.120 ;
  LAYER ME2 ;
  RECT 418.560 0.000 419.680 1.120 ;
  LAYER ME1 ;
  RECT 418.560 0.000 419.680 1.120 ;
 END
END DO24
PIN DI24
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER ME3 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER ME2 ;
  RECT 409.880 0.000 411.000 1.120 ;
  LAYER ME1 ;
  RECT 409.880 0.000 411.000 1.120 ;
 END
END DI24
PIN DO23
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER ME3 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER ME2 ;
  RECT 404.920 0.000 406.040 1.120 ;
  LAYER ME1 ;
  RECT 404.920 0.000 406.040 1.120 ;
 END
END DO23
PIN DI23
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 396.860 0.000 397.980 1.120 ;
  LAYER ME3 ;
  RECT 396.860 0.000 397.980 1.120 ;
  LAYER ME2 ;
  RECT 396.860 0.000 397.980 1.120 ;
  LAYER ME1 ;
  RECT 396.860 0.000 397.980 1.120 ;
 END
END DI23
PIN DO22
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 391.900 0.000 393.020 1.120 ;
  LAYER ME3 ;
  RECT 391.900 0.000 393.020 1.120 ;
  LAYER ME2 ;
  RECT 391.900 0.000 393.020 1.120 ;
  LAYER ME1 ;
  RECT 391.900 0.000 393.020 1.120 ;
 END
END DO22
PIN DI22
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER ME3 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER ME2 ;
  RECT 383.220 0.000 384.340 1.120 ;
  LAYER ME1 ;
  RECT 383.220 0.000 384.340 1.120 ;
 END
END DI22
PIN DO21
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER ME3 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER ME2 ;
  RECT 375.160 0.000 376.280 1.120 ;
  LAYER ME1 ;
  RECT 375.160 0.000 376.280 1.120 ;
 END
END DO21
PIN DI21
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER ME3 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER ME2 ;
  RECT 367.100 0.000 368.220 1.120 ;
  LAYER ME1 ;
  RECT 367.100 0.000 368.220 1.120 ;
 END
END DI21
PIN DO20
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME3 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME2 ;
  RECT 362.140 0.000 363.260 1.120 ;
  LAYER ME1 ;
  RECT 362.140 0.000 363.260 1.120 ;
 END
END DO20
PIN DI20
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 353.460 0.000 354.580 1.120 ;
  LAYER ME3 ;
  RECT 353.460 0.000 354.580 1.120 ;
  LAYER ME2 ;
  RECT 353.460 0.000 354.580 1.120 ;
  LAYER ME1 ;
  RECT 353.460 0.000 354.580 1.120 ;
 END
END DI20
PIN DO19
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME3 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME2 ;
  RECT 348.500 0.000 349.620 1.120 ;
  LAYER ME1 ;
  RECT 348.500 0.000 349.620 1.120 ;
 END
END DO19
PIN DI19
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER ME3 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER ME2 ;
  RECT 340.440 0.000 341.560 1.120 ;
  LAYER ME1 ;
  RECT 340.440 0.000 341.560 1.120 ;
 END
END DI19
PIN DO18
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME3 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME2 ;
  RECT 335.480 0.000 336.600 1.120 ;
  LAYER ME1 ;
  RECT 335.480 0.000 336.600 1.120 ;
 END
END DO18
PIN DI18
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER ME3 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER ME2 ;
  RECT 326.800 0.000 327.920 1.120 ;
  LAYER ME1 ;
  RECT 326.800 0.000 327.920 1.120 ;
 END
END DI18
PIN DO17
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER ME3 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER ME2 ;
  RECT 318.740 0.000 319.860 1.120 ;
  LAYER ME1 ;
  RECT 318.740 0.000 319.860 1.120 ;
 END
END DO17
PIN DI17
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 310.060 0.000 311.180 1.120 ;
  LAYER ME3 ;
  RECT 310.060 0.000 311.180 1.120 ;
  LAYER ME2 ;
  RECT 310.060 0.000 311.180 1.120 ;
  LAYER ME1 ;
  RECT 310.060 0.000 311.180 1.120 ;
 END
END DI17
PIN DO16
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER ME3 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER ME2 ;
  RECT 305.100 0.000 306.220 1.120 ;
  LAYER ME1 ;
  RECT 305.100 0.000 306.220 1.120 ;
 END
END DO16
PIN DI16
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 297.040 0.000 298.160 1.120 ;
  LAYER ME3 ;
  RECT 297.040 0.000 298.160 1.120 ;
  LAYER ME2 ;
  RECT 297.040 0.000 298.160 1.120 ;
  LAYER ME1 ;
  RECT 297.040 0.000 298.160 1.120 ;
 END
END DI16
PIN A1
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 291.460 0.000 292.580 1.120 ;
  LAYER ME3 ;
  RECT 291.460 0.000 292.580 1.120 ;
  LAYER ME2 ;
  RECT 291.460 0.000 292.580 1.120 ;
  LAYER ME1 ;
  RECT 291.460 0.000 292.580 1.120 ;
 END
END A1
PIN WEB
  DIRECTION INPUT ;
  CAPACITANCE 0.011 ;
 PORT
  LAYER ME4 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME3 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME2 ;
  RECT 289.600 0.000 290.720 1.120 ;
  LAYER ME1 ;
  RECT 289.600 0.000 290.720 1.120 ;
 END
END WEB
PIN OE
  DIRECTION INPUT ;
  CAPACITANCE 0.033 ;
 PORT
  LAYER ME4 ;
  RECT 284.640 0.000 285.760 1.120 ;
  LAYER ME3 ;
  RECT 284.640 0.000 285.760 1.120 ;
  LAYER ME2 ;
  RECT 284.640 0.000 285.760 1.120 ;
  LAYER ME1 ;
  RECT 284.640 0.000 285.760 1.120 ;
 END
END OE
PIN CS
  DIRECTION INPUT ;
  CAPACITANCE 0.123 ;
 PORT
  LAYER ME4 ;
  RECT 282.780 0.000 283.900 1.120 ;
  LAYER ME3 ;
  RECT 282.780 0.000 283.900 1.120 ;
  LAYER ME2 ;
  RECT 282.780 0.000 283.900 1.120 ;
  LAYER ME1 ;
  RECT 282.780 0.000 283.900 1.120 ;
 END
END CS
PIN A2
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 261.080 0.000 262.200 1.120 ;
  LAYER ME3 ;
  RECT 261.080 0.000 262.200 1.120 ;
  LAYER ME2 ;
  RECT 261.080 0.000 262.200 1.120 ;
  LAYER ME1 ;
  RECT 261.080 0.000 262.200 1.120 ;
 END
END A2
PIN CK
  DIRECTION INPUT ;
  CAPACITANCE 0.063 ;
 PORT
  LAYER ME4 ;
  RECT 257.980 0.000 259.100 1.120 ;
  LAYER ME3 ;
  RECT 257.980 0.000 259.100 1.120 ;
  LAYER ME2 ;
  RECT 257.980 0.000 259.100 1.120 ;
  LAYER ME1 ;
  RECT 257.980 0.000 259.100 1.120 ;
 END
END CK
PIN A0
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 256.120 0.000 257.240 1.120 ;
  LAYER ME3 ;
  RECT 256.120 0.000 257.240 1.120 ;
  LAYER ME2 ;
  RECT 256.120 0.000 257.240 1.120 ;
  LAYER ME1 ;
  RECT 256.120 0.000 257.240 1.120 ;
 END
END A0
PIN A3
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME3 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME2 ;
  RECT 251.780 0.000 252.900 1.120 ;
  LAYER ME1 ;
  RECT 251.780 0.000 252.900 1.120 ;
 END
END A3
PIN A4
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME3 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME2 ;
  RECT 244.340 0.000 245.460 1.120 ;
  LAYER ME1 ;
  RECT 244.340 0.000 245.460 1.120 ;
 END
END A4
PIN A5
  DIRECTION INPUT ;
  CAPACITANCE 0.027 ;
 PORT
  LAYER ME4 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME3 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME2 ;
  RECT 241.240 0.000 242.360 1.120 ;
  LAYER ME1 ;
  RECT 241.240 0.000 242.360 1.120 ;
 END
END A5
PIN DO15
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME3 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME2 ;
  RECT 233.180 0.000 234.300 1.120 ;
  LAYER ME1 ;
  RECT 233.180 0.000 234.300 1.120 ;
 END
END DO15
PIN DI15
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME3 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME2 ;
  RECT 224.500 0.000 225.620 1.120 ;
  LAYER ME1 ;
  RECT 224.500 0.000 225.620 1.120 ;
 END
END DI15
PIN DO14
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME3 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME2 ;
  RECT 219.540 0.000 220.660 1.120 ;
  LAYER ME1 ;
  RECT 219.540 0.000 220.660 1.120 ;
 END
END DO14
PIN DI14
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME3 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME2 ;
  RECT 211.480 0.000 212.600 1.120 ;
  LAYER ME1 ;
  RECT 211.480 0.000 212.600 1.120 ;
 END
END DI14
PIN DO13
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME3 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME2 ;
  RECT 202.800 0.000 203.920 1.120 ;
  LAYER ME1 ;
  RECT 202.800 0.000 203.920 1.120 ;
 END
END DO13
PIN DI13
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME3 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME2 ;
  RECT 194.740 0.000 195.860 1.120 ;
  LAYER ME1 ;
  RECT 194.740 0.000 195.860 1.120 ;
 END
END DI13
PIN DO12
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME3 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME2 ;
  RECT 189.780 0.000 190.900 1.120 ;
  LAYER ME1 ;
  RECT 189.780 0.000 190.900 1.120 ;
 END
END DO12
PIN DI12
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME3 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME2 ;
  RECT 181.100 0.000 182.220 1.120 ;
  LAYER ME1 ;
  RECT 181.100 0.000 182.220 1.120 ;
 END
END DI12
PIN DO11
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME3 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME2 ;
  RECT 176.140 0.000 177.260 1.120 ;
  LAYER ME1 ;
  RECT 176.140 0.000 177.260 1.120 ;
 END
END DO11
PIN DI11
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME3 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME2 ;
  RECT 168.080 0.000 169.200 1.120 ;
  LAYER ME1 ;
  RECT 168.080 0.000 169.200 1.120 ;
 END
END DI11
PIN DO10
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME3 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME2 ;
  RECT 163.120 0.000 164.240 1.120 ;
  LAYER ME1 ;
  RECT 163.120 0.000 164.240 1.120 ;
 END
END DO10
PIN DI10
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME3 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME2 ;
  RECT 154.440 0.000 155.560 1.120 ;
  LAYER ME1 ;
  RECT 154.440 0.000 155.560 1.120 ;
 END
END DI10
PIN DO9
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME3 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME2 ;
  RECT 146.380 0.000 147.500 1.120 ;
  LAYER ME1 ;
  RECT 146.380 0.000 147.500 1.120 ;
 END
END DO9
PIN DI9
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME3 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME2 ;
  RECT 137.700 0.000 138.820 1.120 ;
  LAYER ME1 ;
  RECT 137.700 0.000 138.820 1.120 ;
 END
END DI9
PIN DO8
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME3 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME2 ;
  RECT 133.360 0.000 134.480 1.120 ;
  LAYER ME1 ;
  RECT 133.360 0.000 134.480 1.120 ;
 END
END DO8
PIN DI8
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME3 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME2 ;
  RECT 124.680 0.000 125.800 1.120 ;
  LAYER ME1 ;
  RECT 124.680 0.000 125.800 1.120 ;
 END
END DI8
PIN DO7
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME3 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME2 ;
  RECT 119.720 0.000 120.840 1.120 ;
  LAYER ME1 ;
  RECT 119.720 0.000 120.840 1.120 ;
 END
END DO7
PIN DI7
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME3 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME2 ;
  RECT 111.660 0.000 112.780 1.120 ;
  LAYER ME1 ;
  RECT 111.660 0.000 112.780 1.120 ;
 END
END DI7
PIN DO6
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME3 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME2 ;
  RECT 106.700 0.000 107.820 1.120 ;
  LAYER ME1 ;
  RECT 106.700 0.000 107.820 1.120 ;
 END
END DO6
PIN DI6
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME3 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME2 ;
  RECT 98.020 0.000 99.140 1.120 ;
  LAYER ME1 ;
  RECT 98.020 0.000 99.140 1.120 ;
 END
END DI6
PIN DO5
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME3 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME2 ;
  RECT 89.960 0.000 91.080 1.120 ;
  LAYER ME1 ;
  RECT 89.960 0.000 91.080 1.120 ;
 END
END DO5
PIN DI5
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME3 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME2 ;
  RECT 81.280 0.000 82.400 1.120 ;
  LAYER ME1 ;
  RECT 81.280 0.000 82.400 1.120 ;
 END
END DI5
PIN DO4
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME3 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME2 ;
  RECT 76.320 0.000 77.440 1.120 ;
  LAYER ME1 ;
  RECT 76.320 0.000 77.440 1.120 ;
 END
END DO4
PIN DI4
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME3 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME2 ;
  RECT 68.260 0.000 69.380 1.120 ;
  LAYER ME1 ;
  RECT 68.260 0.000 69.380 1.120 ;
 END
END DI4
PIN DO3
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME3 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME2 ;
  RECT 63.300 0.000 64.420 1.120 ;
  LAYER ME1 ;
  RECT 63.300 0.000 64.420 1.120 ;
 END
END DO3
PIN DI3
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME3 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME2 ;
  RECT 54.620 0.000 55.740 1.120 ;
  LAYER ME1 ;
  RECT 54.620 0.000 55.740 1.120 ;
 END
END DI3
PIN DO2
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME3 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME2 ;
  RECT 50.280 0.000 51.400 1.120 ;
  LAYER ME1 ;
  RECT 50.280 0.000 51.400 1.120 ;
 END
END DO2
PIN DI2
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME3 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME2 ;
  RECT 41.600 0.000 42.720 1.120 ;
  LAYER ME1 ;
  RECT 41.600 0.000 42.720 1.120 ;
 END
END DI2
PIN DO1
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME3 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME2 ;
  RECT 33.540 0.000 34.660 1.120 ;
  LAYER ME1 ;
  RECT 33.540 0.000 34.660 1.120 ;
 END
END DO1
PIN DI1
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME3 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME2 ;
  RECT 24.860 0.000 25.980 1.120 ;
  LAYER ME1 ;
  RECT 24.860 0.000 25.980 1.120 ;
 END
END DI1
PIN DO0
  DIRECTION OUTPUT ;
  CAPACITANCE 0.031 ;
 PORT
  LAYER ME4 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME3 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME2 ;
  RECT 19.900 0.000 21.020 1.120 ;
  LAYER ME1 ;
  RECT 19.900 0.000 21.020 1.120 ;
 END
END DO0
PIN DI0
  DIRECTION INPUT ;
  CAPACITANCE 0.012 ;
 PORT
  LAYER ME4 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME3 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME2 ;
  RECT 11.840 0.000 12.960 1.120 ;
  LAYER ME1 ;
  RECT 11.840 0.000 12.960 1.120 ;
 END
END DI0
OBS
  LAYER ME1 SPACING 0.280 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER ME2 SPACING 0.320 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER ME3 SPACING 0.320 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER ME4 SPACING 0.600 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER VI1 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER VI2 ;
  RECT 0.000 0.140 531.960 156.800 ;
  LAYER VI3 ;
  RECT 0.000 0.140 531.960 156.800 ;
END
END SRAM_64X32
END LIBRARY



