module PATTERN(
    // Output signals
    clk,
    rst_n,
    cg_en,
    in_valid,
    T,
    in_data,
    w_Q,
    w_K,
    w_V,

    // Input signals
    out_valid,
    out_data
);

output reg clk;
output reg rst_n;
output reg cg_en;
output reg in_valid;
output reg [3:0] T;
output reg signed [7:0] in_data;
output reg signed [7:0] w_Q;
output reg signed [7:0] w_K;
output reg signed [7:0] w_V;

input out_valid;
input signed [63:0] out_data;

//================================================================
// parameters & integer
//================================================================

//================================================================
// Clock
//================================================================
initial clk = 0;
always #(CYCLE/2) clk = ~clk;

//================================================================
// Wire & Reg Declaration
//================================================================


//================================================================
// Task
//================================================================






endmodule